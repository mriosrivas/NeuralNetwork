module log_int(input logic [12:0] in,
	 output logic [15:0] out);
	 	 always_comb
	 	 	 case()
	 	 	 0  : out <= -66019;
	 	 	 1  : out <= -34069;
	 	 	 2  : out <= -31230;
	 	 	 3  : out <= -29569;
	 	 	 4  : out <= -28391;
	 	 	 5  : out <= -27477;
	 	 	 6  : out <= -26730;
	 	 	 7  : out <= -26099;
	 	 	 8  : out <= -25552;
	 	 	 9  : out <= -25069;
	 	 	 10  : out <= -24638;
	 	 	 11  : out <= -24247;
	 	 	 12  : out <= -23891;
	 	 	 13  : out <= -23563;
	 	 	 14  : out <= -23259;
	 	 	 15  : out <= -22977;
	 	 	 16  : out <= -22713;
	 	 	 17  : out <= -22464;
	 	 	 18  : out <= -22230;
	 	 	 19  : out <= -22009;
	 	 	 20  : out <= -21799;
	 	 	 21  : out <= -21599;
	 	 	 22  : out <= -21408;
	 	 	 23  : out <= -21226;
	 	 	 24  : out <= -21052;
	 	 	 25  : out <= -20885;
	 	 	 26  : out <= -20724;
	 	 	 27  : out <= -20569;
	 	 	 28  : out <= -20420;
	 	 	 29  : out <= -20277;
	 	 	 30  : out <= -20138;
	 	 	 31  : out <= -20003;
	 	 	 32  : out <= -19873;
	 	 	 33  : out <= -19747;
	 	 	 34  : out <= -19625;
	 	 	 35  : out <= -19506;
	 	 	 36  : out <= -19391;
	 	 	 37  : out <= -19279;
	 	 	 38  : out <= -19170;
	 	 	 39  : out <= -19063;
	 	 	 40  : out <= -18959;
	 	 	 41  : out <= -18858;
	 	 	 42  : out <= -18760;
	 	 	 43  : out <= -18663;
	 	 	 44  : out <= -18569;
	 	 	 45  : out <= -18477;
	 	 	 46  : out <= -18387;
	 	 	 47  : out <= -18299;
	 	 	 48  : out <= -18213;
	 	 	 49  : out <= -18128;
	 	 	 50  : out <= -18045;
	 	 	 51  : out <= -17964;
	 	 	 52  : out <= -17885;
	 	 	 53  : out <= -17807;
	 	 	 54  : out <= -17730;
	 	 	 55  : out <= -17655;
	 	 	 56  : out <= -17581;
	 	 	 57  : out <= -17509;
	 	 	 58  : out <= -17437;
	 	 	 59  : out <= -17367;
	 	 	 60  : out <= -17299;
	 	 	 61  : out <= -17231;
	 	 	 62  : out <= -17164;
	 	 	 63  : out <= -17099;
	 	 	 64  : out <= -17034;
	 	 	 65  : out <= -16971;
	 	 	 66  : out <= -16908;
	 	 	 67  : out <= -16847;
	 	 	 68  : out <= -16786;
	 	 	 69  : out <= -16726;
	 	 	 70  : out <= -16667;
	 	 	 71  : out <= -16609;
	 	 	 72  : out <= -16552;
	 	 	 73  : out <= -16495;
	 	 	 74  : out <= -16440;
	 	 	 75  : out <= -16385;
	 	 	 76  : out <= -16330;
	 	 	 77  : out <= -16277;
	 	 	 78  : out <= -16224;
	 	 	 79  : out <= -16172;
	 	 	 80  : out <= -16120;
	 	 	 81  : out <= -16069;
	 	 	 82  : out <= -16019;
	 	 	 83  : out <= -15969;
	 	 	 84  : out <= -15920;
	 	 	 85  : out <= -15872;
	 	 	 86  : out <= -15824;
	 	 	 87  : out <= -15777;
	 	 	 88  : out <= -15730;
	 	 	 89  : out <= -15684;
	 	 	 90  : out <= -15638;
	 	 	 91  : out <= -15593;
	 	 	 92  : out <= -15548;
	 	 	 93  : out <= -15504;
	 	 	 94  : out <= -15460;
	 	 	 95  : out <= -15416;
	 	 	 96  : out <= -15374;
	 	 	 97  : out <= -15331;
	 	 	 98  : out <= -15289;
	 	 	 99  : out <= -15247;
	 	 	 100  : out <= -15206;
	 	 	 101  : out <= -15166;
	 	 	 102  : out <= -15125;
	 	 	 103  : out <= -15085;
	 	 	 104  : out <= -15046;
	 	 	 105  : out <= -15006;
	 	 	 106  : out <= -14968;
	 	 	 107  : out <= -14929;
	 	 	 108  : out <= -14891;
	 	 	 109  : out <= -14853;
	 	 	 110  : out <= -14816;
	 	 	 111  : out <= -14779;
	 	 	 112  : out <= -14742;
	 	 	 113  : out <= -14706;
	 	 	 114  : out <= -14670;
	 	 	 115  : out <= -14634;
	 	 	 116  : out <= -14598;
	 	 	 117  : out <= -14563;
	 	 	 118  : out <= -14528;
	 	 	 119  : out <= -14494;
	 	 	 120  : out <= -14460;
	 	 	 121  : out <= -14426;
	 	 	 122  : out <= -14392;
	 	 	 123  : out <= -14358;
	 	 	 124  : out <= -14325;
	 	 	 125  : out <= -14292;
	 	 	 126  : out <= -14260;
	 	 	 127  : out <= -14227;
	 	 	 128  : out <= -14195;
	 	 	 129  : out <= -14163;
	 	 	 130  : out <= -14132;
	 	 	 131  : out <= -14100;
	 	 	 132  : out <= -14069;
	 	 	 133  : out <= -14038;
	 	 	 134  : out <= -14008;
	 	 	 135  : out <= -13977;
	 	 	 136  : out <= -13947;
	 	 	 137  : out <= -13917;
	 	 	 138  : out <= -13887;
	 	 	 139  : out <= -13857;
	 	 	 140  : out <= -13828;
	 	 	 141  : out <= -13799;
	 	 	 142  : out <= -13770;
	 	 	 143  : out <= -13741;
	 	 	 144  : out <= -13713;
	 	 	 145  : out <= -13684;
	 	 	 146  : out <= -13656;
	 	 	 147  : out <= -13628;
	 	 	 148  : out <= -13600;
	 	 	 149  : out <= -13573;
	 	 	 150  : out <= -13546;
	 	 	 151  : out <= -13518;
	 	 	 152  : out <= -13491;
	 	 	 153  : out <= -13464;
	 	 	 154  : out <= -13438;
	 	 	 155  : out <= -13411;
	 	 	 156  : out <= -13385;
	 	 	 157  : out <= -13359;
	 	 	 158  : out <= -13333;
	 	 	 159  : out <= -13307;
	 	 	 160  : out <= -13281;
	 	 	 161  : out <= -13256;
	 	 	 162  : out <= -13230;
	 	 	 163  : out <= -13205;
	 	 	 164  : out <= -13180;
	 	 	 165  : out <= -13155;
	 	 	 166  : out <= -13130;
	 	 	 167  : out <= -13106;
	 	 	 168  : out <= -13081;
	 	 	 169  : out <= -13057;
	 	 	 170  : out <= -13033;
	 	 	 171  : out <= -13009;
	 	 	 172  : out <= -12985;
	 	 	 173  : out <= -12961;
	 	 	 174  : out <= -12938;
	 	 	 175  : out <= -12914;
	 	 	 176  : out <= -12891;
	 	 	 177  : out <= -12868;
	 	 	 178  : out <= -12844;
	 	 	 179  : out <= -12822;
	 	 	 180  : out <= -12799;
	 	 	 181  : out <= -12776;
	 	 	 182  : out <= -12753;
	 	 	 183  : out <= -12731;
	 	 	 184  : out <= -12709;
	 	 	 185  : out <= -12686;
	 	 	 186  : out <= -12664;
	 	 	 187  : out <= -12642;
	 	 	 188  : out <= -12621;
	 	 	 189  : out <= -12599;
	 	 	 190  : out <= -12577;
	 	 	 191  : out <= -12556;
	 	 	 192  : out <= -12534;
	 	 	 193  : out <= -12513;
	 	 	 194  : out <= -12492;
	 	 	 195  : out <= -12471;
	 	 	 196  : out <= -12450;
	 	 	 197  : out <= -12429;
	 	 	 198  : out <= -12408;
	 	 	 199  : out <= -12388;
	 	 	 200  : out <= -12367;
	 	 	 201  : out <= -12347;
	 	 	 202  : out <= -12326;
	 	 	 203  : out <= -12306;
	 	 	 204  : out <= -12286;
	 	 	 205  : out <= -12266;
	 	 	 206  : out <= -12246;
	 	 	 207  : out <= -12226;
	 	 	 208  : out <= -12207;
	 	 	 209  : out <= -12187;
	 	 	 210  : out <= -12167;
	 	 	 211  : out <= -12148;
	 	 	 212  : out <= -12128;
	 	 	 213  : out <= -12109;
	 	 	 214  : out <= -12090;
	 	 	 215  : out <= -12071;
	 	 	 216  : out <= -12052;
	 	 	 217  : out <= -12033;
	 	 	 218  : out <= -12014;
	 	 	 219  : out <= -11995;
	 	 	 220  : out <= -11977;
	 	 	 221  : out <= -11958;
	 	 	 222  : out <= -11940;
	 	 	 223  : out <= -11921;
	 	 	 224  : out <= -11903;
	 	 	 225  : out <= -11885;
	 	 	 226  : out <= -11867;
	 	 	 227  : out <= -11848;
	 	 	 228  : out <= -11830;
	 	 	 229  : out <= -11813;
	 	 	 230  : out <= -11795;
	 	 	 231  : out <= -11777;
	 	 	 232  : out <= -11759;
	 	 	 233  : out <= -11742;
	 	 	 234  : out <= -11724;
	 	 	 235  : out <= -11707;
	 	 	 236  : out <= -11689;
	 	 	 237  : out <= -11672;
	 	 	 238  : out <= -11655;
	 	 	 239  : out <= -11637;
	 	 	 240  : out <= -11620;
	 	 	 241  : out <= -11603;
	 	 	 242  : out <= -11586;
	 	 	 243  : out <= -11569;
	 	 	 244  : out <= -11553;
	 	 	 245  : out <= -11536;
	 	 	 246  : out <= -11519;
	 	 	 247  : out <= -11503;
	 	 	 248  : out <= -11486;
	 	 	 249  : out <= -11470;
	 	 	 250  : out <= -11453;
	 	 	 251  : out <= -11437;
	 	 	 252  : out <= -11421;
	 	 	 253  : out <= -11404;
	 	 	 254  : out <= -11388;
	 	 	 255  : out <= -11372;
	 	 	 256  : out <= -11356;
	 	 	 257  : out <= -11340;
	 	 	 258  : out <= -11324;
	 	 	 259  : out <= -11308;
	 	 	 260  : out <= -11293;
	 	 	 261  : out <= -11277;
	 	 	 262  : out <= -11261;
	 	 	 263  : out <= -11246;
	 	 	 264  : out <= -11230;
	 	 	 265  : out <= -11214;
	 	 	 266  : out <= -11199;
	 	 	 267  : out <= -11184;
	 	 	 268  : out <= -11168;
	 	 	 269  : out <= -11153;
	 	 	 270  : out <= -11138;
	 	 	 271  : out <= -11123;
	 	 	 272  : out <= -11108;
	 	 	 273  : out <= -11093;
	 	 	 274  : out <= -11078;
	 	 	 275  : out <= -11063;
	 	 	 276  : out <= -11048;
	 	 	 277  : out <= -11033;
	 	 	 278  : out <= -11018;
	 	 	 279  : out <= -11004;
	 	 	 280  : out <= -10989;
	 	 	 281  : out <= -10974;
	 	 	 282  : out <= -10960;
	 	 	 283  : out <= -10945;
	 	 	 284  : out <= -10931;
	 	 	 285  : out <= -10916;
	 	 	 286  : out <= -10902;
	 	 	 287  : out <= -10888;
	 	 	 288  : out <= -10874;
	 	 	 289  : out <= -10859;
	 	 	 290  : out <= -10845;
	 	 	 291  : out <= -10831;
	 	 	 292  : out <= -10817;
	 	 	 293  : out <= -10803;
	 	 	 294  : out <= -10789;
	 	 	 295  : out <= -10775;
	 	 	 296  : out <= -10761;
	 	 	 297  : out <= -10748;
	 	 	 298  : out <= -10734;
	 	 	 299  : out <= -10720;
	 	 	 300  : out <= -10706;
	 	 	 301  : out <= -10693;
	 	 	 302  : out <= -10679;
	 	 	 303  : out <= -10666;
	 	 	 304  : out <= -10652;
	 	 	 305  : out <= -10639;
	 	 	 306  : out <= -10625;
	 	 	 307  : out <= -10612;
	 	 	 308  : out <= -10599;
	 	 	 309  : out <= -10585;
	 	 	 310  : out <= -10572;
	 	 	 311  : out <= -10559;
	 	 	 312  : out <= -10546;
	 	 	 313  : out <= -10533;
	 	 	 314  : out <= -10520;
	 	 	 315  : out <= -10507;
	 	 	 316  : out <= -10494;
	 	 	 317  : out <= -10481;
	 	 	 318  : out <= -10468;
	 	 	 319  : out <= -10455;
	 	 	 320  : out <= -10442;
	 	 	 321  : out <= -10429;
	 	 	 322  : out <= -10417;
	 	 	 323  : out <= -10404;
	 	 	 324  : out <= -10391;
	 	 	 325  : out <= -10379;
	 	 	 326  : out <= -10366;
	 	 	 327  : out <= -10353;
	 	 	 328  : out <= -10341;
	 	 	 329  : out <= -10328;
	 	 	 330  : out <= -10316;
	 	 	 331  : out <= -10304;
	 	 	 332  : out <= -10291;
	 	 	 333  : out <= -10279;
	 	 	 334  : out <= -10267;
	 	 	 335  : out <= -10254;
	 	 	 336  : out <= -10242;
	 	 	 337  : out <= -10230;
	 	 	 338  : out <= -10218;
	 	 	 339  : out <= -10206;
	 	 	 340  : out <= -10194;
	 	 	 341  : out <= -10182;
	 	 	 342  : out <= -10170;
	 	 	 343  : out <= -10158;
	 	 	 344  : out <= -10146;
	 	 	 345  : out <= -10134;
	 	 	 346  : out <= -10122;
	 	 	 347  : out <= -10110;
	 	 	 348  : out <= -10098;
	 	 	 349  : out <= -10087;
	 	 	 350  : out <= -10075;
	 	 	 351  : out <= -10063;
	 	 	 352  : out <= -10052;
	 	 	 353  : out <= -10040;
	 	 	 354  : out <= -10028;
	 	 	 355  : out <= -10017;
	 	 	 356  : out <= -10005;
	 	 	 357  : out <= -9994;
	 	 	 358  : out <= -9982;
	 	 	 359  : out <= -9971;
	 	 	 360  : out <= -9960;
	 	 	 361  : out <= -9948;
	 	 	 362  : out <= -9937;
	 	 	 363  : out <= -9926;
	 	 	 364  : out <= -9914;
	 	 	 365  : out <= -9903;
	 	 	 366  : out <= -9892;
	 	 	 367  : out <= -9881;
	 	 	 368  : out <= -9870;
	 	 	 369  : out <= -9858;
	 	 	 370  : out <= -9847;
	 	 	 371  : out <= -9836;
	 	 	 372  : out <= -9825;
	 	 	 373  : out <= -9814;
	 	 	 374  : out <= -9803;
	 	 	 375  : out <= -9792;
	 	 	 376  : out <= -9781;
	 	 	 377  : out <= -9771;
	 	 	 378  : out <= -9760;
	 	 	 379  : out <= -9749;
	 	 	 380  : out <= -9738;
	 	 	 381  : out <= -9727;
	 	 	 382  : out <= -9717;
	 	 	 383  : out <= -9706;
	 	 	 384  : out <= -9695;
	 	 	 385  : out <= -9685;
	 	 	 386  : out <= -9674;
	 	 	 387  : out <= -9663;
	 	 	 388  : out <= -9653;
	 	 	 389  : out <= -9642;
	 	 	 390  : out <= -9632;
	 	 	 391  : out <= -9621;
	 	 	 392  : out <= -9611;
	 	 	 393  : out <= -9600;
	 	 	 394  : out <= -9590;
	 	 	 395  : out <= -9580;
	 	 	 396  : out <= -9569;
	 	 	 397  : out <= -9559;
	 	 	 398  : out <= -9549;
	 	 	 399  : out <= -9538;
	 	 	 400  : out <= -9528;
	 	 	 401  : out <= -9518;
	 	 	 402  : out <= -9508;
	 	 	 403  : out <= -9497;
	 	 	 404  : out <= -9487;
	 	 	 405  : out <= -9477;
	 	 	 406  : out <= -9467;
	 	 	 407  : out <= -9457;
	 	 	 408  : out <= -9447;
	 	 	 409  : out <= -9437;
	 	 	 410  : out <= -9427;
	 	 	 411  : out <= -9417;
	 	 	 412  : out <= -9407;
	 	 	 413  : out <= -9397;
	 	 	 414  : out <= -9387;
	 	 	 415  : out <= -9377;
	 	 	 416  : out <= -9367;
	 	 	 417  : out <= -9358;
	 	 	 418  : out <= -9348;
	 	 	 419  : out <= -9338;
	 	 	 420  : out <= -9328;
	 	 	 421  : out <= -9318;
	 	 	 422  : out <= -9309;
	 	 	 423  : out <= -9299;
	 	 	 424  : out <= -9289;
	 	 	 425  : out <= -9280;
	 	 	 426  : out <= -9270;
	 	 	 427  : out <= -9260;
	 	 	 428  : out <= -9251;
	 	 	 429  : out <= -9241;
	 	 	 430  : out <= -9232;
	 	 	 431  : out <= -9222;
	 	 	 432  : out <= -9213;
	 	 	 433  : out <= -9203;
	 	 	 434  : out <= -9194;
	 	 	 435  : out <= -9184;
	 	 	 436  : out <= -9175;
	 	 	 437  : out <= -9166;
	 	 	 438  : out <= -9156;
	 	 	 439  : out <= -9147;
	 	 	 440  : out <= -9138;
	 	 	 441  : out <= -9128;
	 	 	 442  : out <= -9119;
	 	 	 443  : out <= -9110;
	 	 	 444  : out <= -9101;
	 	 	 445  : out <= -9091;
	 	 	 446  : out <= -9082;
	 	 	 447  : out <= -9073;
	 	 	 448  : out <= -9064;
	 	 	 449  : out <= -9055;
	 	 	 450  : out <= -9046;
	 	 	 451  : out <= -9036;
	 	 	 452  : out <= -9027;
	 	 	 453  : out <= -9018;
	 	 	 454  : out <= -9009;
	 	 	 455  : out <= -9000;
	 	 	 456  : out <= -8991;
	 	 	 457  : out <= -8982;
	 	 	 458  : out <= -8973;
	 	 	 459  : out <= -8964;
	 	 	 460  : out <= -8956;
	 	 	 461  : out <= -8947;
	 	 	 462  : out <= -8938;
	 	 	 463  : out <= -8929;
	 	 	 464  : out <= -8920;
	 	 	 465  : out <= -8911;
	 	 	 466  : out <= -8902;
	 	 	 467  : out <= -8894;
	 	 	 468  : out <= -8885;
	 	 	 469  : out <= -8876;
	 	 	 470  : out <= -8867;
	 	 	 471  : out <= -8859;
	 	 	 472  : out <= -8850;
	 	 	 473  : out <= -8841;
	 	 	 474  : out <= -8833;
	 	 	 475  : out <= -8824;
	 	 	 476  : out <= -8816;
	 	 	 477  : out <= -8807;
	 	 	 478  : out <= -8798;
	 	 	 479  : out <= -8790;
	 	 	 480  : out <= -8781;
	 	 	 481  : out <= -8773;
	 	 	 482  : out <= -8764;
	 	 	 483  : out <= -8756;
	 	 	 484  : out <= -8747;
	 	 	 485  : out <= -8739;
	 	 	 486  : out <= -8730;
	 	 	 487  : out <= -8722;
	 	 	 488  : out <= -8714;
	 	 	 489  : out <= -8705;
	 	 	 490  : out <= -8697;
	 	 	 491  : out <= -8688;
	 	 	 492  : out <= -8680;
	 	 	 493  : out <= -8672;
	 	 	 494  : out <= -8663;
	 	 	 495  : out <= -8655;
	 	 	 496  : out <= -8647;
	 	 	 497  : out <= -8639;
	 	 	 498  : out <= -8630;
	 	 	 499  : out <= -8622;
	 	 	 500  : out <= -8614;
	 	 	 501  : out <= -8606;
	 	 	 502  : out <= -8598;
	 	 	 503  : out <= -8590;
	 	 	 504  : out <= -8581;
	 	 	 505  : out <= -8573;
	 	 	 506  : out <= -8565;
	 	 	 507  : out <= -8557;
	 	 	 508  : out <= -8549;
	 	 	 509  : out <= -8541;
	 	 	 510  : out <= -8533;
	 	 	 511  : out <= -8525;
	 	 	 512  : out <= -8517;
	 	 	 513  : out <= -8509;
	 	 	 514  : out <= -8501;
	 	 	 515  : out <= -8493;
	 	 	 516  : out <= -8485;
	 	 	 517  : out <= -8477;
	 	 	 518  : out <= -8469;
	 	 	 519  : out <= -8461;
	 	 	 520  : out <= -8453;
	 	 	 521  : out <= -8446;
	 	 	 522  : out <= -8438;
	 	 	 523  : out <= -8430;
	 	 	 524  : out <= -8422;
	 	 	 525  : out <= -8414;
	 	 	 526  : out <= -8406;
	 	 	 527  : out <= -8399;
	 	 	 528  : out <= -8391;
	 	 	 529  : out <= -8383;
	 	 	 530  : out <= -8375;
	 	 	 531  : out <= -8368;
	 	 	 532  : out <= -8360;
	 	 	 533  : out <= -8352;
	 	 	 534  : out <= -8345;
	 	 	 535  : out <= -8337;
	 	 	 536  : out <= -8329;
	 	 	 537  : out <= -8322;
	 	 	 538  : out <= -8314;
	 	 	 539  : out <= -8306;
	 	 	 540  : out <= -8299;
	 	 	 541  : out <= -8291;
	 	 	 542  : out <= -8284;
	 	 	 543  : out <= -8276;
	 	 	 544  : out <= -8269;
	 	 	 545  : out <= -8261;
	 	 	 546  : out <= -8254;
	 	 	 547  : out <= -8246;
	 	 	 548  : out <= -8239;
	 	 	 549  : out <= -8231;
	 	 	 550  : out <= -8224;
	 	 	 551  : out <= -8216;
	 	 	 552  : out <= -8209;
	 	 	 553  : out <= -8201;
	 	 	 554  : out <= -8194;
	 	 	 555  : out <= -8187;
	 	 	 556  : out <= -8179;
	 	 	 557  : out <= -8172;
	 	 	 558  : out <= -8164;
	 	 	 559  : out <= -8157;
	 	 	 560  : out <= -8150;
	 	 	 561  : out <= -8143;
	 	 	 562  : out <= -8135;
	 	 	 563  : out <= -8128;
	 	 	 564  : out <= -8121;
	 	 	 565  : out <= -8113;
	 	 	 566  : out <= -8106;
	 	 	 567  : out <= -8099;
	 	 	 568  : out <= -8092;
	 	 	 569  : out <= -8085;
	 	 	 570  : out <= -8077;
	 	 	 571  : out <= -8070;
	 	 	 572  : out <= -8063;
	 	 	 573  : out <= -8056;
	 	 	 574  : out <= -8049;
	 	 	 575  : out <= -8042;
	 	 	 576  : out <= -8034;
	 	 	 577  : out <= -8027;
	 	 	 578  : out <= -8020;
	 	 	 579  : out <= -8013;
	 	 	 580  : out <= -8006;
	 	 	 581  : out <= -7999;
	 	 	 582  : out <= -7992;
	 	 	 583  : out <= -7985;
	 	 	 584  : out <= -7978;
	 	 	 585  : out <= -7971;
	 	 	 586  : out <= -7964;
	 	 	 587  : out <= -7957;
	 	 	 588  : out <= -7950;
	 	 	 589  : out <= -7943;
	 	 	 590  : out <= -7936;
	 	 	 591  : out <= -7929;
	 	 	 592  : out <= -7922;
	 	 	 593  : out <= -7915;
	 	 	 594  : out <= -7908;
	 	 	 595  : out <= -7902;
	 	 	 596  : out <= -7895;
	 	 	 597  : out <= -7888;
	 	 	 598  : out <= -7881;
	 	 	 599  : out <= -7874;
	 	 	 600  : out <= -7867;
	 	 	 601  : out <= -7860;
	 	 	 602  : out <= -7854;
	 	 	 603  : out <= -7847;
	 	 	 604  : out <= -7840;
	 	 	 605  : out <= -7833;
	 	 	 606  : out <= -7826;
	 	 	 607  : out <= -7820;
	 	 	 608  : out <= -7813;
	 	 	 609  : out <= -7806;
	 	 	 610  : out <= -7800;
	 	 	 611  : out <= -7793;
	 	 	 612  : out <= -7786;
	 	 	 613  : out <= -7779;
	 	 	 614  : out <= -7773;
	 	 	 615  : out <= -7766;
	 	 	 616  : out <= -7759;
	 	 	 617  : out <= -7753;
	 	 	 618  : out <= -7746;
	 	 	 619  : out <= -7740;
	 	 	 620  : out <= -7733;
	 	 	 621  : out <= -7726;
	 	 	 622  : out <= -7720;
	 	 	 623  : out <= -7713;
	 	 	 624  : out <= -7707;
	 	 	 625  : out <= -7700;
	 	 	 626  : out <= -7693;
	 	 	 627  : out <= -7687;
	 	 	 628  : out <= -7680;
	 	 	 629  : out <= -7674;
	 	 	 630  : out <= -7667;
	 	 	 631  : out <= -7661;
	 	 	 632  : out <= -7654;
	 	 	 633  : out <= -7648;
	 	 	 634  : out <= -7641;
	 	 	 635  : out <= -7635;
	 	 	 636  : out <= -7629;
	 	 	 637  : out <= -7622;
	 	 	 638  : out <= -7616;
	 	 	 639  : out <= -7609;
	 	 	 640  : out <= -7603;
	 	 	 641  : out <= -7597;
	 	 	 642  : out <= -7590;
	 	 	 643  : out <= -7584;
	 	 	 644  : out <= -7577;
	 	 	 645  : out <= -7571;
	 	 	 646  : out <= -7565;
	 	 	 647  : out <= -7558;
	 	 	 648  : out <= -7552;
	 	 	 649  : out <= -7546;
	 	 	 650  : out <= -7539;
	 	 	 651  : out <= -7533;
	 	 	 652  : out <= -7527;
	 	 	 653  : out <= -7521;
	 	 	 654  : out <= -7514;
	 	 	 655  : out <= -7508;
	 	 	 656  : out <= -7502;
	 	 	 657  : out <= -7496;
	 	 	 658  : out <= -7489;
	 	 	 659  : out <= -7483;
	 	 	 660  : out <= -7477;
	 	 	 661  : out <= -7471;
	 	 	 662  : out <= -7464;
	 	 	 663  : out <= -7458;
	 	 	 664  : out <= -7452;
	 	 	 665  : out <= -7446;
	 	 	 666  : out <= -7440;
	 	 	 667  : out <= -7434;
	 	 	 668  : out <= -7428;
	 	 	 669  : out <= -7421;
	 	 	 670  : out <= -7415;
	 	 	 671  : out <= -7409;
	 	 	 672  : out <= -7403;
	 	 	 673  : out <= -7397;
	 	 	 674  : out <= -7391;
	 	 	 675  : out <= -7385;
	 	 	 676  : out <= -7379;
	 	 	 677  : out <= -7373;
	 	 	 678  : out <= -7367;
	 	 	 679  : out <= -7361;
	 	 	 680  : out <= -7355;
	 	 	 681  : out <= -7349;
	 	 	 682  : out <= -7343;
	 	 	 683  : out <= -7337;
	 	 	 684  : out <= -7331;
	 	 	 685  : out <= -7325;
	 	 	 686  : out <= -7319;
	 	 	 687  : out <= -7313;
	 	 	 688  : out <= -7307;
	 	 	 689  : out <= -7301;
	 	 	 690  : out <= -7295;
	 	 	 691  : out <= -7289;
	 	 	 692  : out <= -7283;
	 	 	 693  : out <= -7277;
	 	 	 694  : out <= -7271;
	 	 	 695  : out <= -7265;
	 	 	 696  : out <= -7259;
	 	 	 697  : out <= -7253;
	 	 	 698  : out <= -7248;
	 	 	 699  : out <= -7242;
	 	 	 700  : out <= -7236;
	 	 	 701  : out <= -7230;
	 	 	 702  : out <= -7224;
	 	 	 703  : out <= -7218;
	 	 	 704  : out <= -7213;
	 	 	 705  : out <= -7207;
	 	 	 706  : out <= -7201;
	 	 	 707  : out <= -7195;
	 	 	 708  : out <= -7189;
	 	 	 709  : out <= -7184;
	 	 	 710  : out <= -7178;
	 	 	 711  : out <= -7172;
	 	 	 712  : out <= -7166;
	 	 	 713  : out <= -7160;
	 	 	 714  : out <= -7155;
	 	 	 715  : out <= -7149;
	 	 	 716  : out <= -7143;
	 	 	 717  : out <= -7138;
	 	 	 718  : out <= -7132;
	 	 	 719  : out <= -7126;
	 	 	 720  : out <= -7120;
	 	 	 721  : out <= -7115;
	 	 	 722  : out <= -7109;
	 	 	 723  : out <= -7103;
	 	 	 724  : out <= -7098;
	 	 	 725  : out <= -7092;
	 	 	 726  : out <= -7086;
	 	 	 727  : out <= -7081;
	 	 	 728  : out <= -7075;
	 	 	 729  : out <= -7070;
	 	 	 730  : out <= -7064;
	 	 	 731  : out <= -7058;
	 	 	 732  : out <= -7053;
	 	 	 733  : out <= -7047;
	 	 	 734  : out <= -7042;
	 	 	 735  : out <= -7036;
	 	 	 736  : out <= -7030;
	 	 	 737  : out <= -7025;
	 	 	 738  : out <= -7019;
	 	 	 739  : out <= -7014;
	 	 	 740  : out <= -7008;
	 	 	 741  : out <= -7003;
	 	 	 742  : out <= -6997;
	 	 	 743  : out <= -6992;
	 	 	 744  : out <= -6986;
	 	 	 745  : out <= -6981;
	 	 	 746  : out <= -6975;
	 	 	 747  : out <= -6970;
	 	 	 748  : out <= -6964;
	 	 	 749  : out <= -6959;
	 	 	 750  : out <= -6953;
	 	 	 751  : out <= -6948;
	 	 	 752  : out <= -6942;
	 	 	 753  : out <= -6937;
	 	 	 754  : out <= -6931;
	 	 	 755  : out <= -6926;
	 	 	 756  : out <= -6921;
	 	 	 757  : out <= -6915;
	 	 	 758  : out <= -6910;
	 	 	 759  : out <= -6904;
	 	 	 760  : out <= -6899;
	 	 	 761  : out <= -6894;
	 	 	 762  : out <= -6888;
	 	 	 763  : out <= -6883;
	 	 	 764  : out <= -6877;
	 	 	 765  : out <= -6872;
	 	 	 766  : out <= -6867;
	 	 	 767  : out <= -6861;
	 	 	 768  : out <= -6856;
	 	 	 769  : out <= -6851;
	 	 	 770  : out <= -6845;
	 	 	 771  : out <= -6840;
	 	 	 772  : out <= -6835;
	 	 	 773  : out <= -6830;
	 	 	 774  : out <= -6824;
	 	 	 775  : out <= -6819;
	 	 	 776  : out <= -6814;
	 	 	 777  : out <= -6808;
	 	 	 778  : out <= -6803;
	 	 	 779  : out <= -6798;
	 	 	 780  : out <= -6793;
	 	 	 781  : out <= -6787;
	 	 	 782  : out <= -6782;
	 	 	 783  : out <= -6777;
	 	 	 784  : out <= -6772;
	 	 	 785  : out <= -6766;
	 	 	 786  : out <= -6761;
	 	 	 787  : out <= -6756;
	 	 	 788  : out <= -6751;
	 	 	 789  : out <= -6746;
	 	 	 790  : out <= -6740;
	 	 	 791  : out <= -6735;
	 	 	 792  : out <= -6730;
	 	 	 793  : out <= -6725;
	 	 	 794  : out <= -6720;
	 	 	 795  : out <= -6715;
	 	 	 796  : out <= -6709;
	 	 	 797  : out <= -6704;
	 	 	 798  : out <= -6699;
	 	 	 799  : out <= -6694;
	 	 	 800  : out <= -6689;
	 	 	 801  : out <= -6684;
	 	 	 802  : out <= -6679;
	 	 	 803  : out <= -6674;
	 	 	 804  : out <= -6668;
	 	 	 805  : out <= -6663;
	 	 	 806  : out <= -6658;
	 	 	 807  : out <= -6653;
	 	 	 808  : out <= -6648;
	 	 	 809  : out <= -6643;
	 	 	 810  : out <= -6638;
	 	 	 811  : out <= -6633;
	 	 	 812  : out <= -6628;
	 	 	 813  : out <= -6623;
	 	 	 814  : out <= -6618;
	 	 	 815  : out <= -6613;
	 	 	 816  : out <= -6608;
	 	 	 817  : out <= -6603;
	 	 	 818  : out <= -6598;
	 	 	 819  : out <= -6593;
	 	 	 820  : out <= -6588;
	 	 	 821  : out <= -6583;
	 	 	 822  : out <= -6578;
	 	 	 823  : out <= -6573;
	 	 	 824  : out <= -6568;
	 	 	 825  : out <= -6563;
	 	 	 826  : out <= -6558;
	 	 	 827  : out <= -6553;
	 	 	 828  : out <= -6548;
	 	 	 829  : out <= -6543;
	 	 	 830  : out <= -6538;
	 	 	 831  : out <= -6533;
	 	 	 832  : out <= -6528;
	 	 	 833  : out <= -6523;
	 	 	 834  : out <= -6518;
	 	 	 835  : out <= -6514;
	 	 	 836  : out <= -6509;
	 	 	 837  : out <= -6504;
	 	 	 838  : out <= -6499;
	 	 	 839  : out <= -6494;
	 	 	 840  : out <= -6489;
	 	 	 841  : out <= -6484;
	 	 	 842  : out <= -6479;
	 	 	 843  : out <= -6474;
	 	 	 844  : out <= -6470;
	 	 	 845  : out <= -6465;
	 	 	 846  : out <= -6460;
	 	 	 847  : out <= -6455;
	 	 	 848  : out <= -6450;
	 	 	 849  : out <= -6445;
	 	 	 850  : out <= -6441;
	 	 	 851  : out <= -6436;
	 	 	 852  : out <= -6431;
	 	 	 853  : out <= -6426;
	 	 	 854  : out <= -6421;
	 	 	 855  : out <= -6417;
	 	 	 856  : out <= -6412;
	 	 	 857  : out <= -6407;
	 	 	 858  : out <= -6402;
	 	 	 859  : out <= -6397;
	 	 	 860  : out <= -6393;
	 	 	 861  : out <= -6388;
	 	 	 862  : out <= -6383;
	 	 	 863  : out <= -6378;
	 	 	 864  : out <= -6374;
	 	 	 865  : out <= -6369;
	 	 	 866  : out <= -6364;
	 	 	 867  : out <= -6359;
	 	 	 868  : out <= -6355;
	 	 	 869  : out <= -6350;
	 	 	 870  : out <= -6345;
	 	 	 871  : out <= -6341;
	 	 	 872  : out <= -6336;
	 	 	 873  : out <= -6331;
	 	 	 874  : out <= -6327;
	 	 	 875  : out <= -6322;
	 	 	 876  : out <= -6317;
	 	 	 877  : out <= -6312;
	 	 	 878  : out <= -6308;
	 	 	 879  : out <= -6303;
	 	 	 880  : out <= -6299;
	 	 	 881  : out <= -6294;
	 	 	 882  : out <= -6289;
	 	 	 883  : out <= -6285;
	 	 	 884  : out <= -6280;
	 	 	 885  : out <= -6275;
	 	 	 886  : out <= -6271;
	 	 	 887  : out <= -6266;
	 	 	 888  : out <= -6261;
	 	 	 889  : out <= -6257;
	 	 	 890  : out <= -6252;
	 	 	 891  : out <= -6248;
	 	 	 892  : out <= -6243;
	 	 	 893  : out <= -6238;
	 	 	 894  : out <= -6234;
	 	 	 895  : out <= -6229;
	 	 	 896  : out <= -6225;
	 	 	 897  : out <= -6220;
	 	 	 898  : out <= -6216;
	 	 	 899  : out <= -6211;
	 	 	 900  : out <= -6206;
	 	 	 901  : out <= -6202;
	 	 	 902  : out <= -6197;
	 	 	 903  : out <= -6193;
	 	 	 904  : out <= -6188;
	 	 	 905  : out <= -6184;
	 	 	 906  : out <= -6179;
	 	 	 907  : out <= -6175;
	 	 	 908  : out <= -6170;
	 	 	 909  : out <= -6166;
	 	 	 910  : out <= -6161;
	 	 	 911  : out <= -6157;
	 	 	 912  : out <= -6152;
	 	 	 913  : out <= -6148;
	 	 	 914  : out <= -6143;
	 	 	 915  : out <= -6139;
	 	 	 916  : out <= -6134;
	 	 	 917  : out <= -6130;
	 	 	 918  : out <= -6125;
	 	 	 919  : out <= -6121;
	 	 	 920  : out <= -6116;
	 	 	 921  : out <= -6112;
	 	 	 922  : out <= -6108;
	 	 	 923  : out <= -6103;
	 	 	 924  : out <= -6099;
	 	 	 925  : out <= -6094;
	 	 	 926  : out <= -6090;
	 	 	 927  : out <= -6085;
	 	 	 928  : out <= -6081;
	 	 	 929  : out <= -6077;
	 	 	 930  : out <= -6072;
	 	 	 931  : out <= -6068;
	 	 	 932  : out <= -6063;
	 	 	 933  : out <= -6059;
	 	 	 934  : out <= -6055;
	 	 	 935  : out <= -6050;
	 	 	 936  : out <= -6046;
	 	 	 937  : out <= -6041;
	 	 	 938  : out <= -6037;
	 	 	 939  : out <= -6033;
	 	 	 940  : out <= -6028;
	 	 	 941  : out <= -6024;
	 	 	 942  : out <= -6020;
	 	 	 943  : out <= -6015;
	 	 	 944  : out <= -6011;
	 	 	 945  : out <= -6007;
	 	 	 946  : out <= -6002;
	 	 	 947  : out <= -5998;
	 	 	 948  : out <= -5994;
	 	 	 949  : out <= -5989;
	 	 	 950  : out <= -5985;
	 	 	 951  : out <= -5981;
	 	 	 952  : out <= -5976;
	 	 	 953  : out <= -5972;
	 	 	 954  : out <= -5968;
	 	 	 955  : out <= -5964;
	 	 	 956  : out <= -5959;
	 	 	 957  : out <= -5955;
	 	 	 958  : out <= -5951;
	 	 	 959  : out <= -5946;
	 	 	 960  : out <= -5942;
	 	 	 961  : out <= -5938;
	 	 	 962  : out <= -5934;
	 	 	 963  : out <= -5929;
	 	 	 964  : out <= -5925;
	 	 	 965  : out <= -5921;
	 	 	 966  : out <= -5917;
	 	 	 967  : out <= -5912;
	 	 	 968  : out <= -5908;
	 	 	 969  : out <= -5904;
	 	 	 970  : out <= -5900;
	 	 	 971  : out <= -5895;
	 	 	 972  : out <= -5891;
	 	 	 973  : out <= -5887;
	 	 	 974  : out <= -5883;
	 	 	 975  : out <= -5879;
	 	 	 976  : out <= -5874;
	 	 	 977  : out <= -5870;
	 	 	 978  : out <= -5866;
	 	 	 979  : out <= -5862;
	 	 	 980  : out <= -5858;
	 	 	 981  : out <= -5853;
	 	 	 982  : out <= -5849;
	 	 	 983  : out <= -5845;
	 	 	 984  : out <= -5841;
	 	 	 985  : out <= -5837;
	 	 	 986  : out <= -5833;
	 	 	 987  : out <= -5829;
	 	 	 988  : out <= -5824;
	 	 	 989  : out <= -5820;
	 	 	 990  : out <= -5816;
	 	 	 991  : out <= -5812;
	 	 	 992  : out <= -5808;
	 	 	 993  : out <= -5804;
	 	 	 994  : out <= -5800;
	 	 	 995  : out <= -5795;
	 	 	 996  : out <= -5791;
	 	 	 997  : out <= -5787;
	 	 	 998  : out <= -5783;
	 	 	 999  : out <= -5779;
	 	 	 1000  : out <= -5775;
	 	 	 1001  : out <= -5771;
	 	 	 1002  : out <= -5767;
	 	 	 1003  : out <= -5763;
	 	 	 1004  : out <= -5759;
	 	 	 1005  : out <= -5754;
	 	 	 1006  : out <= -5750;
	 	 	 1007  : out <= -5746;
	 	 	 1008  : out <= -5742;
	 	 	 1009  : out <= -5738;
	 	 	 1010  : out <= -5734;
	 	 	 1011  : out <= -5730;
	 	 	 1012  : out <= -5726;
	 	 	 1013  : out <= -5722;
	 	 	 1014  : out <= -5718;
	 	 	 1015  : out <= -5714;
	 	 	 1016  : out <= -5710;
	 	 	 1017  : out <= -5706;
	 	 	 1018  : out <= -5702;
	 	 	 1019  : out <= -5698;
	 	 	 1020  : out <= -5694;
	 	 	 1021  : out <= -5690;
	 	 	 1022  : out <= -5686;
	 	 	 1023  : out <= -5682;
	 	 	 1024  : out <= -5678;
	 	 	 1025  : out <= -5674;
	 	 	 1026  : out <= -5670;
	 	 	 1027  : out <= -5666;
	 	 	 1028  : out <= -5662;
	 	 	 1029  : out <= -5658;
	 	 	 1030  : out <= -5654;
	 	 	 1031  : out <= -5650;
	 	 	 1032  : out <= -5646;
	 	 	 1033  : out <= -5642;
	 	 	 1034  : out <= -5638;
	 	 	 1035  : out <= -5634;
	 	 	 1036  : out <= -5630;
	 	 	 1037  : out <= -5626;
	 	 	 1038  : out <= -5622;
	 	 	 1039  : out <= -5618;
	 	 	 1040  : out <= -5614;
	 	 	 1041  : out <= -5610;
	 	 	 1042  : out <= -5606;
	 	 	 1043  : out <= -5602;
	 	 	 1044  : out <= -5599;
	 	 	 1045  : out <= -5595;
	 	 	 1046  : out <= -5591;
	 	 	 1047  : out <= -5587;
	 	 	 1048  : out <= -5583;
	 	 	 1049  : out <= -5579;
	 	 	 1050  : out <= -5575;
	 	 	 1051  : out <= -5571;
	 	 	 1052  : out <= -5567;
	 	 	 1053  : out <= -5563;
	 	 	 1054  : out <= -5559;
	 	 	 1055  : out <= -5556;
	 	 	 1056  : out <= -5552;
	 	 	 1057  : out <= -5548;
	 	 	 1058  : out <= -5544;
	 	 	 1059  : out <= -5540;
	 	 	 1060  : out <= -5536;
	 	 	 1061  : out <= -5532;
	 	 	 1062  : out <= -5529;
	 	 	 1063  : out <= -5525;
	 	 	 1064  : out <= -5521;
	 	 	 1065  : out <= -5517;
	 	 	 1066  : out <= -5513;
	 	 	 1067  : out <= -5509;
	 	 	 1068  : out <= -5505;
	 	 	 1069  : out <= -5502;
	 	 	 1070  : out <= -5498;
	 	 	 1071  : out <= -5494;
	 	 	 1072  : out <= -5490;
	 	 	 1073  : out <= -5486;
	 	 	 1074  : out <= -5482;
	 	 	 1075  : out <= -5479;
	 	 	 1076  : out <= -5475;
	 	 	 1077  : out <= -5471;
	 	 	 1078  : out <= -5467;
	 	 	 1079  : out <= -5463;
	 	 	 1080  : out <= -5460;
	 	 	 1081  : out <= -5456;
	 	 	 1082  : out <= -5452;
	 	 	 1083  : out <= -5448;
	 	 	 1084  : out <= -5445;
	 	 	 1085  : out <= -5441;
	 	 	 1086  : out <= -5437;
	 	 	 1087  : out <= -5433;
	 	 	 1088  : out <= -5429;
	 	 	 1089  : out <= -5426;
	 	 	 1090  : out <= -5422;
	 	 	 1091  : out <= -5418;
	 	 	 1092  : out <= -5414;
	 	 	 1093  : out <= -5411;
	 	 	 1094  : out <= -5407;
	 	 	 1095  : out <= -5403;
	 	 	 1096  : out <= -5399;
	 	 	 1097  : out <= -5396;
	 	 	 1098  : out <= -5392;
	 	 	 1099  : out <= -5388;
	 	 	 1100  : out <= -5385;
	 	 	 1101  : out <= -5381;
	 	 	 1102  : out <= -5377;
	 	 	 1103  : out <= -5373;
	 	 	 1104  : out <= -5370;
	 	 	 1105  : out <= -5366;
	 	 	 1106  : out <= -5362;
	 	 	 1107  : out <= -5359;
	 	 	 1108  : out <= -5355;
	 	 	 1109  : out <= -5351;
	 	 	 1110  : out <= -5347;
	 	 	 1111  : out <= -5344;
	 	 	 1112  : out <= -5340;
	 	 	 1113  : out <= -5336;
	 	 	 1114  : out <= -5333;
	 	 	 1115  : out <= -5329;
	 	 	 1116  : out <= -5325;
	 	 	 1117  : out <= -5322;
	 	 	 1118  : out <= -5318;
	 	 	 1119  : out <= -5314;
	 	 	 1120  : out <= -5311;
	 	 	 1121  : out <= -5307;
	 	 	 1122  : out <= -5303;
	 	 	 1123  : out <= -5300;
	 	 	 1124  : out <= -5296;
	 	 	 1125  : out <= -5292;
	 	 	 1126  : out <= -5289;
	 	 	 1127  : out <= -5285;
	 	 	 1128  : out <= -5282;
	 	 	 1129  : out <= -5278;
	 	 	 1130  : out <= -5274;
	 	 	 1131  : out <= -5271;
	 	 	 1132  : out <= -5267;
	 	 	 1133  : out <= -5263;
	 	 	 1134  : out <= -5260;
	 	 	 1135  : out <= -5256;
	 	 	 1136  : out <= -5253;
	 	 	 1137  : out <= -5249;
	 	 	 1138  : out <= -5245;
	 	 	 1139  : out <= -5242;
	 	 	 1140  : out <= -5238;
	 	 	 1141  : out <= -5235;
	 	 	 1142  : out <= -5231;
	 	 	 1143  : out <= -5227;
	 	 	 1144  : out <= -5224;
	 	 	 1145  : out <= -5220;
	 	 	 1146  : out <= -5217;
	 	 	 1147  : out <= -5213;
	 	 	 1148  : out <= -5210;
	 	 	 1149  : out <= -5206;
	 	 	 1150  : out <= -5202;
	 	 	 1151  : out <= -5199;
	 	 	 1152  : out <= -5195;
	 	 	 1153  : out <= -5192;
	 	 	 1154  : out <= -5188;
	 	 	 1155  : out <= -5185;
	 	 	 1156  : out <= -5181;
	 	 	 1157  : out <= -5178;
	 	 	 1158  : out <= -5174;
	 	 	 1159  : out <= -5171;
	 	 	 1160  : out <= -5167;
	 	 	 1161  : out <= -5163;
	 	 	 1162  : out <= -5160;
	 	 	 1163  : out <= -5156;
	 	 	 1164  : out <= -5153;
	 	 	 1165  : out <= -5149;
	 	 	 1166  : out <= -5146;
	 	 	 1167  : out <= -5142;
	 	 	 1168  : out <= -5139;
	 	 	 1169  : out <= -5135;
	 	 	 1170  : out <= -5132;
	 	 	 1171  : out <= -5128;
	 	 	 1172  : out <= -5125;
	 	 	 1173  : out <= -5121;
	 	 	 1174  : out <= -5118;
	 	 	 1175  : out <= -5114;
	 	 	 1176  : out <= -5111;
	 	 	 1177  : out <= -5107;
	 	 	 1178  : out <= -5104;
	 	 	 1179  : out <= -5100;
	 	 	 1180  : out <= -5097;
	 	 	 1181  : out <= -5093;
	 	 	 1182  : out <= -5090;
	 	 	 1183  : out <= -5087;
	 	 	 1184  : out <= -5083;
	 	 	 1185  : out <= -5080;
	 	 	 1186  : out <= -5076;
	 	 	 1187  : out <= -5073;
	 	 	 1188  : out <= -5069;
	 	 	 1189  : out <= -5066;
	 	 	 1190  : out <= -5062;
	 	 	 1191  : out <= -5059;
	 	 	 1192  : out <= -5056;
	 	 	 1193  : out <= -5052;
	 	 	 1194  : out <= -5049;
	 	 	 1195  : out <= -5045;
	 	 	 1196  : out <= -5042;
	 	 	 1197  : out <= -5038;
	 	 	 1198  : out <= -5035;
	 	 	 1199  : out <= -5032;
	 	 	 1200  : out <= -5028;
	 	 	 1201  : out <= -5025;
	 	 	 1202  : out <= -5021;
	 	 	 1203  : out <= -5018;
	 	 	 1204  : out <= -5014;
	 	 	 1205  : out <= -5011;
	 	 	 1206  : out <= -5008;
	 	 	 1207  : out <= -5004;
	 	 	 1208  : out <= -5001;
	 	 	 1209  : out <= -4998;
	 	 	 1210  : out <= -4994;
	 	 	 1211  : out <= -4991;
	 	 	 1212  : out <= -4987;
	 	 	 1213  : out <= -4984;
	 	 	 1214  : out <= -4981;
	 	 	 1215  : out <= -4977;
	 	 	 1216  : out <= -4974;
	 	 	 1217  : out <= -4970;
	 	 	 1218  : out <= -4967;
	 	 	 1219  : out <= -4964;
	 	 	 1220  : out <= -4960;
	 	 	 1221  : out <= -4957;
	 	 	 1222  : out <= -4954;
	 	 	 1223  : out <= -4950;
	 	 	 1224  : out <= -4947;
	 	 	 1225  : out <= -4944;
	 	 	 1226  : out <= -4940;
	 	 	 1227  : out <= -4937;
	 	 	 1228  : out <= -4934;
	 	 	 1229  : out <= -4930;
	 	 	 1230  : out <= -4927;
	 	 	 1231  : out <= -4924;
	 	 	 1232  : out <= -4920;
	 	 	 1233  : out <= -4917;
	 	 	 1234  : out <= -4914;
	 	 	 1235  : out <= -4910;
	 	 	 1236  : out <= -4907;
	 	 	 1237  : out <= -4904;
	 	 	 1238  : out <= -4900;
	 	 	 1239  : out <= -4897;
	 	 	 1240  : out <= -4894;
	 	 	 1241  : out <= -4891;
	 	 	 1242  : out <= -4887;
	 	 	 1243  : out <= -4884;
	 	 	 1244  : out <= -4881;
	 	 	 1245  : out <= -4877;
	 	 	 1246  : out <= -4874;
	 	 	 1247  : out <= -4871;
	 	 	 1248  : out <= -4867;
	 	 	 1249  : out <= -4864;
	 	 	 1250  : out <= -4861;
	 	 	 1251  : out <= -4858;
	 	 	 1252  : out <= -4854;
	 	 	 1253  : out <= -4851;
	 	 	 1254  : out <= -4848;
	 	 	 1255  : out <= -4845;
	 	 	 1256  : out <= -4841;
	 	 	 1257  : out <= -4838;
	 	 	 1258  : out <= -4835;
	 	 	 1259  : out <= -4832;
	 	 	 1260  : out <= -4828;
	 	 	 1261  : out <= -4825;
	 	 	 1262  : out <= -4822;
	 	 	 1263  : out <= -4819;
	 	 	 1264  : out <= -4815;
	 	 	 1265  : out <= -4812;
	 	 	 1266  : out <= -4809;
	 	 	 1267  : out <= -4806;
	 	 	 1268  : out <= -4802;
	 	 	 1269  : out <= -4799;
	 	 	 1270  : out <= -4796;
	 	 	 1271  : out <= -4793;
	 	 	 1272  : out <= -4789;
	 	 	 1273  : out <= -4786;
	 	 	 1274  : out <= -4783;
	 	 	 1275  : out <= -4780;
	 	 	 1276  : out <= -4777;
	 	 	 1277  : out <= -4773;
	 	 	 1278  : out <= -4770;
	 	 	 1279  : out <= -4767;
	 	 	 1280  : out <= -4764;
	 	 	 1281  : out <= -4761;
	 	 	 1282  : out <= -4757;
	 	 	 1283  : out <= -4754;
	 	 	 1284  : out <= -4751;
	 	 	 1285  : out <= -4748;
	 	 	 1286  : out <= -4745;
	 	 	 1287  : out <= -4741;
	 	 	 1288  : out <= -4738;
	 	 	 1289  : out <= -4735;
	 	 	 1290  : out <= -4732;
	 	 	 1291  : out <= -4729;
	 	 	 1292  : out <= -4726;
	 	 	 1293  : out <= -4722;
	 	 	 1294  : out <= -4719;
	 	 	 1295  : out <= -4716;
	 	 	 1296  : out <= -4713;
	 	 	 1297  : out <= -4710;
	 	 	 1298  : out <= -4707;
	 	 	 1299  : out <= -4703;
	 	 	 1300  : out <= -4700;
	 	 	 1301  : out <= -4697;
	 	 	 1302  : out <= -4694;
	 	 	 1303  : out <= -4691;
	 	 	 1304  : out <= -4688;
	 	 	 1305  : out <= -4685;
	 	 	 1306  : out <= -4681;
	 	 	 1307  : out <= -4678;
	 	 	 1308  : out <= -4675;
	 	 	 1309  : out <= -4672;
	 	 	 1310  : out <= -4669;
	 	 	 1311  : out <= -4666;
	 	 	 1312  : out <= -4663;
	 	 	 1313  : out <= -4660;
	 	 	 1314  : out <= -4656;
	 	 	 1315  : out <= -4653;
	 	 	 1316  : out <= -4650;
	 	 	 1317  : out <= -4647;
	 	 	 1318  : out <= -4644;
	 	 	 1319  : out <= -4641;
	 	 	 1320  : out <= -4638;
	 	 	 1321  : out <= -4635;
	 	 	 1322  : out <= -4632;
	 	 	 1323  : out <= -4628;
	 	 	 1324  : out <= -4625;
	 	 	 1325  : out <= -4622;
	 	 	 1326  : out <= -4619;
	 	 	 1327  : out <= -4616;
	 	 	 1328  : out <= -4613;
	 	 	 1329  : out <= -4610;
	 	 	 1330  : out <= -4607;
	 	 	 1331  : out <= -4604;
	 	 	 1332  : out <= -4601;
	 	 	 1333  : out <= -4598;
	 	 	 1334  : out <= -4595;
	 	 	 1335  : out <= -4591;
	 	 	 1336  : out <= -4588;
	 	 	 1337  : out <= -4585;
	 	 	 1338  : out <= -4582;
	 	 	 1339  : out <= -4579;
	 	 	 1340  : out <= -4576;
	 	 	 1341  : out <= -4573;
	 	 	 1342  : out <= -4570;
	 	 	 1343  : out <= -4567;
	 	 	 1344  : out <= -4564;
	 	 	 1345  : out <= -4561;
	 	 	 1346  : out <= -4558;
	 	 	 1347  : out <= -4555;
	 	 	 1348  : out <= -4552;
	 	 	 1349  : out <= -4549;
	 	 	 1350  : out <= -4546;
	 	 	 1351  : out <= -4543;
	 	 	 1352  : out <= -4540;
	 	 	 1353  : out <= -4537;
	 	 	 1354  : out <= -4534;
	 	 	 1355  : out <= -4531;
	 	 	 1356  : out <= -4528;
	 	 	 1357  : out <= -4524;
	 	 	 1358  : out <= -4521;
	 	 	 1359  : out <= -4518;
	 	 	 1360  : out <= -4515;
	 	 	 1361  : out <= -4512;
	 	 	 1362  : out <= -4509;
	 	 	 1363  : out <= -4506;
	 	 	 1364  : out <= -4503;
	 	 	 1365  : out <= -4500;
	 	 	 1366  : out <= -4497;
	 	 	 1367  : out <= -4494;
	 	 	 1368  : out <= -4491;
	 	 	 1369  : out <= -4488;
	 	 	 1370  : out <= -4485;
	 	 	 1371  : out <= -4482;
	 	 	 1372  : out <= -4479;
	 	 	 1373  : out <= -4476;
	 	 	 1374  : out <= -4473;
	 	 	 1375  : out <= -4471;
	 	 	 1376  : out <= -4468;
	 	 	 1377  : out <= -4465;
	 	 	 1378  : out <= -4462;
	 	 	 1379  : out <= -4459;
	 	 	 1380  : out <= -4456;
	 	 	 1381  : out <= -4453;
	 	 	 1382  : out <= -4450;
	 	 	 1383  : out <= -4447;
	 	 	 1384  : out <= -4444;
	 	 	 1385  : out <= -4441;
	 	 	 1386  : out <= -4438;
	 	 	 1387  : out <= -4435;
	 	 	 1388  : out <= -4432;
	 	 	 1389  : out <= -4429;
	 	 	 1390  : out <= -4426;
	 	 	 1391  : out <= -4423;
	 	 	 1392  : out <= -4420;
	 	 	 1393  : out <= -4417;
	 	 	 1394  : out <= -4414;
	 	 	 1395  : out <= -4411;
	 	 	 1396  : out <= -4408;
	 	 	 1397  : out <= -4406;
	 	 	 1398  : out <= -4403;
	 	 	 1399  : out <= -4400;
	 	 	 1400  : out <= -4397;
	 	 	 1401  : out <= -4394;
	 	 	 1402  : out <= -4391;
	 	 	 1403  : out <= -4388;
	 	 	 1404  : out <= -4385;
	 	 	 1405  : out <= -4382;
	 	 	 1406  : out <= -4379;
	 	 	 1407  : out <= -4376;
	 	 	 1408  : out <= -4373;
	 	 	 1409  : out <= -4370;
	 	 	 1410  : out <= -4368;
	 	 	 1411  : out <= -4365;
	 	 	 1412  : out <= -4362;
	 	 	 1413  : out <= -4359;
	 	 	 1414  : out <= -4356;
	 	 	 1415  : out <= -4353;
	 	 	 1416  : out <= -4350;
	 	 	 1417  : out <= -4347;
	 	 	 1418  : out <= -4344;
	 	 	 1419  : out <= -4341;
	 	 	 1420  : out <= -4339;
	 	 	 1421  : out <= -4336;
	 	 	 1422  : out <= -4333;
	 	 	 1423  : out <= -4330;
	 	 	 1424  : out <= -4327;
	 	 	 1425  : out <= -4324;
	 	 	 1426  : out <= -4321;
	 	 	 1427  : out <= -4318;
	 	 	 1428  : out <= -4316;
	 	 	 1429  : out <= -4313;
	 	 	 1430  : out <= -4310;
	 	 	 1431  : out <= -4307;
	 	 	 1432  : out <= -4304;
	 	 	 1433  : out <= -4301;
	 	 	 1434  : out <= -4298;
	 	 	 1435  : out <= -4296;
	 	 	 1436  : out <= -4293;
	 	 	 1437  : out <= -4290;
	 	 	 1438  : out <= -4287;
	 	 	 1439  : out <= -4284;
	 	 	 1440  : out <= -4281;
	 	 	 1441  : out <= -4278;
	 	 	 1442  : out <= -4276;
	 	 	 1443  : out <= -4273;
	 	 	 1444  : out <= -4270;
	 	 	 1445  : out <= -4267;
	 	 	 1446  : out <= -4264;
	 	 	 1447  : out <= -4261;
	 	 	 1448  : out <= -4259;
	 	 	 1449  : out <= -4256;
	 	 	 1450  : out <= -4253;
	 	 	 1451  : out <= -4250;
	 	 	 1452  : out <= -4247;
	 	 	 1453  : out <= -4245;
	 	 	 1454  : out <= -4242;
	 	 	 1455  : out <= -4239;
	 	 	 1456  : out <= -4236;
	 	 	 1457  : out <= -4233;
	 	 	 1458  : out <= -4230;
	 	 	 1459  : out <= -4228;
	 	 	 1460  : out <= -4225;
	 	 	 1461  : out <= -4222;
	 	 	 1462  : out <= -4219;
	 	 	 1463  : out <= -4216;
	 	 	 1464  : out <= -4214;
	 	 	 1465  : out <= -4211;
	 	 	 1466  : out <= -4208;
	 	 	 1467  : out <= -4205;
	 	 	 1468  : out <= -4202;
	 	 	 1469  : out <= -4200;
	 	 	 1470  : out <= -4197;
	 	 	 1471  : out <= -4194;
	 	 	 1472  : out <= -4191;
	 	 	 1473  : out <= -4189;
	 	 	 1474  : out <= -4186;
	 	 	 1475  : out <= -4183;
	 	 	 1476  : out <= -4180;
	 	 	 1477  : out <= -4177;
	 	 	 1478  : out <= -4175;
	 	 	 1479  : out <= -4172;
	 	 	 1480  : out <= -4169;
	 	 	 1481  : out <= -4166;
	 	 	 1482  : out <= -4164;
	 	 	 1483  : out <= -4161;
	 	 	 1484  : out <= -4158;
	 	 	 1485  : out <= -4155;
	 	 	 1486  : out <= -4153;
	 	 	 1487  : out <= -4150;
	 	 	 1488  : out <= -4147;
	 	 	 1489  : out <= -4144;
	 	 	 1490  : out <= -4142;
	 	 	 1491  : out <= -4139;
	 	 	 1492  : out <= -4136;
	 	 	 1493  : out <= -4133;
	 	 	 1494  : out <= -4131;
	 	 	 1495  : out <= -4128;
	 	 	 1496  : out <= -4125;
	 	 	 1497  : out <= -4122;
	 	 	 1498  : out <= -4120;
	 	 	 1499  : out <= -4117;
	 	 	 1500  : out <= -4114;
	 	 	 1501  : out <= -4111;
	 	 	 1502  : out <= -4109;
	 	 	 1503  : out <= -4106;
	 	 	 1504  : out <= -4103;
	 	 	 1505  : out <= -4100;
	 	 	 1506  : out <= -4098;
	 	 	 1507  : out <= -4095;
	 	 	 1508  : out <= -4092;
	 	 	 1509  : out <= -4090;
	 	 	 1510  : out <= -4087;
	 	 	 1511  : out <= -4084;
	 	 	 1512  : out <= -4081;
	 	 	 1513  : out <= -4079;
	 	 	 1514  : out <= -4076;
	 	 	 1515  : out <= -4073;
	 	 	 1516  : out <= -4071;
	 	 	 1517  : out <= -4068;
	 	 	 1518  : out <= -4065;
	 	 	 1519  : out <= -4063;
	 	 	 1520  : out <= -4060;
	 	 	 1521  : out <= -4057;
	 	 	 1522  : out <= -4054;
	 	 	 1523  : out <= -4052;
	 	 	 1524  : out <= -4049;
	 	 	 1525  : out <= -4046;
	 	 	 1526  : out <= -4044;
	 	 	 1527  : out <= -4041;
	 	 	 1528  : out <= -4038;
	 	 	 1529  : out <= -4036;
	 	 	 1530  : out <= -4033;
	 	 	 1531  : out <= -4030;
	 	 	 1532  : out <= -4028;
	 	 	 1533  : out <= -4025;
	 	 	 1534  : out <= -4022;
	 	 	 1535  : out <= -4020;
	 	 	 1536  : out <= -4017;
	 	 	 1537  : out <= -4014;
	 	 	 1538  : out <= -4012;
	 	 	 1539  : out <= -4009;
	 	 	 1540  : out <= -4006;
	 	 	 1541  : out <= -4004;
	 	 	 1542  : out <= -4001;
	 	 	 1543  : out <= -3998;
	 	 	 1544  : out <= -3996;
	 	 	 1545  : out <= -3993;
	 	 	 1546  : out <= -3990;
	 	 	 1547  : out <= -3988;
	 	 	 1548  : out <= -3985;
	 	 	 1549  : out <= -3982;
	 	 	 1550  : out <= -3980;
	 	 	 1551  : out <= -3977;
	 	 	 1552  : out <= -3975;
	 	 	 1553  : out <= -3972;
	 	 	 1554  : out <= -3969;
	 	 	 1555  : out <= -3967;
	 	 	 1556  : out <= -3964;
	 	 	 1557  : out <= -3961;
	 	 	 1558  : out <= -3959;
	 	 	 1559  : out <= -3956;
	 	 	 1560  : out <= -3953;
	 	 	 1561  : out <= -3951;
	 	 	 1562  : out <= -3948;
	 	 	 1563  : out <= -3946;
	 	 	 1564  : out <= -3943;
	 	 	 1565  : out <= -3940;
	 	 	 1566  : out <= -3938;
	 	 	 1567  : out <= -3935;
	 	 	 1568  : out <= -3933;
	 	 	 1569  : out <= -3930;
	 	 	 1570  : out <= -3927;
	 	 	 1571  : out <= -3925;
	 	 	 1572  : out <= -3922;
	 	 	 1573  : out <= -3919;
	 	 	 1574  : out <= -3917;
	 	 	 1575  : out <= -3914;
	 	 	 1576  : out <= -3912;
	 	 	 1577  : out <= -3909;
	 	 	 1578  : out <= -3906;
	 	 	 1579  : out <= -3904;
	 	 	 1580  : out <= -3901;
	 	 	 1581  : out <= -3899;
	 	 	 1582  : out <= -3896;
	 	 	 1583  : out <= -3894;
	 	 	 1584  : out <= -3891;
	 	 	 1585  : out <= -3888;
	 	 	 1586  : out <= -3886;
	 	 	 1587  : out <= -3883;
	 	 	 1588  : out <= -3881;
	 	 	 1589  : out <= -3878;
	 	 	 1590  : out <= -3875;
	 	 	 1591  : out <= -3873;
	 	 	 1592  : out <= -3870;
	 	 	 1593  : out <= -3868;
	 	 	 1594  : out <= -3865;
	 	 	 1595  : out <= -3863;
	 	 	 1596  : out <= -3860;
	 	 	 1597  : out <= -3857;
	 	 	 1598  : out <= -3855;
	 	 	 1599  : out <= -3852;
	 	 	 1600  : out <= -3850;
	 	 	 1601  : out <= -3847;
	 	 	 1602  : out <= -3845;
	 	 	 1603  : out <= -3842;
	 	 	 1604  : out <= -3840;
	 	 	 1605  : out <= -3837;
	 	 	 1606  : out <= -3834;
	 	 	 1607  : out <= -3832;
	 	 	 1608  : out <= -3829;
	 	 	 1609  : out <= -3827;
	 	 	 1610  : out <= -3824;
	 	 	 1611  : out <= -3822;
	 	 	 1612  : out <= -3819;
	 	 	 1613  : out <= -3817;
	 	 	 1614  : out <= -3814;
	 	 	 1615  : out <= -3812;
	 	 	 1616  : out <= -3809;
	 	 	 1617  : out <= -3806;
	 	 	 1618  : out <= -3804;
	 	 	 1619  : out <= -3801;
	 	 	 1620  : out <= -3799;
	 	 	 1621  : out <= -3796;
	 	 	 1622  : out <= -3794;
	 	 	 1623  : out <= -3791;
	 	 	 1624  : out <= -3789;
	 	 	 1625  : out <= -3786;
	 	 	 1626  : out <= -3784;
	 	 	 1627  : out <= -3781;
	 	 	 1628  : out <= -3779;
	 	 	 1629  : out <= -3776;
	 	 	 1630  : out <= -3774;
	 	 	 1631  : out <= -3771;
	 	 	 1632  : out <= -3769;
	 	 	 1633  : out <= -3766;
	 	 	 1634  : out <= -3764;
	 	 	 1635  : out <= -3761;
	 	 	 1636  : out <= -3759;
	 	 	 1637  : out <= -3756;
	 	 	 1638  : out <= -3754;
	 	 	 1639  : out <= -3751;
	 	 	 1640  : out <= -3749;
	 	 	 1641  : out <= -3746;
	 	 	 1642  : out <= -3744;
	 	 	 1643  : out <= -3741;
	 	 	 1644  : out <= -3739;
	 	 	 1645  : out <= -3736;
	 	 	 1646  : out <= -3734;
	 	 	 1647  : out <= -3731;
	 	 	 1648  : out <= -3729;
	 	 	 1649  : out <= -3726;
	 	 	 1650  : out <= -3724;
	 	 	 1651  : out <= -3721;
	 	 	 1652  : out <= -3719;
	 	 	 1653  : out <= -3716;
	 	 	 1654  : out <= -3714;
	 	 	 1655  : out <= -3711;
	 	 	 1656  : out <= -3709;
	 	 	 1657  : out <= -3706;
	 	 	 1658  : out <= -3704;
	 	 	 1659  : out <= -3701;
	 	 	 1660  : out <= -3699;
	 	 	 1661  : out <= -3697;
	 	 	 1662  : out <= -3694;
	 	 	 1663  : out <= -3692;
	 	 	 1664  : out <= -3689;
	 	 	 1665  : out <= -3687;
	 	 	 1666  : out <= -3684;
	 	 	 1667  : out <= -3682;
	 	 	 1668  : out <= -3679;
	 	 	 1669  : out <= -3677;
	 	 	 1670  : out <= -3674;
	 	 	 1671  : out <= -3672;
	 	 	 1672  : out <= -3669;
	 	 	 1673  : out <= -3667;
	 	 	 1674  : out <= -3665;
	 	 	 1675  : out <= -3662;
	 	 	 1676  : out <= -3660;
	 	 	 1677  : out <= -3657;
	 	 	 1678  : out <= -3655;
	 	 	 1679  : out <= -3652;
	 	 	 1680  : out <= -3650;
	 	 	 1681  : out <= -3647;
	 	 	 1682  : out <= -3645;
	 	 	 1683  : out <= -3643;
	 	 	 1684  : out <= -3640;
	 	 	 1685  : out <= -3638;
	 	 	 1686  : out <= -3635;
	 	 	 1687  : out <= -3633;
	 	 	 1688  : out <= -3630;
	 	 	 1689  : out <= -3628;
	 	 	 1690  : out <= -3626;
	 	 	 1691  : out <= -3623;
	 	 	 1692  : out <= -3621;
	 	 	 1693  : out <= -3618;
	 	 	 1694  : out <= -3616;
	 	 	 1695  : out <= -3614;
	 	 	 1696  : out <= -3611;
	 	 	 1697  : out <= -3609;
	 	 	 1698  : out <= -3606;
	 	 	 1699  : out <= -3604;
	 	 	 1700  : out <= -3601;
	 	 	 1701  : out <= -3599;
	 	 	 1702  : out <= -3597;
	 	 	 1703  : out <= -3594;
	 	 	 1704  : out <= -3592;
	 	 	 1705  : out <= -3589;
	 	 	 1706  : out <= -3587;
	 	 	 1707  : out <= -3585;
	 	 	 1708  : out <= -3582;
	 	 	 1709  : out <= -3580;
	 	 	 1710  : out <= -3577;
	 	 	 1711  : out <= -3575;
	 	 	 1712  : out <= -3573;
	 	 	 1713  : out <= -3570;
	 	 	 1714  : out <= -3568;
	 	 	 1715  : out <= -3565;
	 	 	 1716  : out <= -3563;
	 	 	 1717  : out <= -3561;
	 	 	 1718  : out <= -3558;
	 	 	 1719  : out <= -3556;
	 	 	 1720  : out <= -3554;
	 	 	 1721  : out <= -3551;
	 	 	 1722  : out <= -3549;
	 	 	 1723  : out <= -3546;
	 	 	 1724  : out <= -3544;
	 	 	 1725  : out <= -3542;
	 	 	 1726  : out <= -3539;
	 	 	 1727  : out <= -3537;
	 	 	 1728  : out <= -3535;
	 	 	 1729  : out <= -3532;
	 	 	 1730  : out <= -3530;
	 	 	 1731  : out <= -3527;
	 	 	 1732  : out <= -3525;
	 	 	 1733  : out <= -3523;
	 	 	 1734  : out <= -3520;
	 	 	 1735  : out <= -3518;
	 	 	 1736  : out <= -3516;
	 	 	 1737  : out <= -3513;
	 	 	 1738  : out <= -3511;
	 	 	 1739  : out <= -3509;
	 	 	 1740  : out <= -3506;
	 	 	 1741  : out <= -3504;
	 	 	 1742  : out <= -3501;
	 	 	 1743  : out <= -3499;
	 	 	 1744  : out <= -3497;
	 	 	 1745  : out <= -3494;
	 	 	 1746  : out <= -3492;
	 	 	 1747  : out <= -3490;
	 	 	 1748  : out <= -3487;
	 	 	 1749  : out <= -3485;
	 	 	 1750  : out <= -3483;
	 	 	 1751  : out <= -3480;
	 	 	 1752  : out <= -3478;
	 	 	 1753  : out <= -3476;
	 	 	 1754  : out <= -3473;
	 	 	 1755  : out <= -3471;
	 	 	 1756  : out <= -3469;
	 	 	 1757  : out <= -3466;
	 	 	 1758  : out <= -3464;
	 	 	 1759  : out <= -3462;
	 	 	 1760  : out <= -3459;
	 	 	 1761  : out <= -3457;
	 	 	 1762  : out <= -3455;
	 	 	 1763  : out <= -3452;
	 	 	 1764  : out <= -3450;
	 	 	 1765  : out <= -3448;
	 	 	 1766  : out <= -3445;
	 	 	 1767  : out <= -3443;
	 	 	 1768  : out <= -3441;
	 	 	 1769  : out <= -3438;
	 	 	 1770  : out <= -3436;
	 	 	 1771  : out <= -3434;
	 	 	 1772  : out <= -3432;
	 	 	 1773  : out <= -3429;
	 	 	 1774  : out <= -3427;
	 	 	 1775  : out <= -3425;
	 	 	 1776  : out <= -3422;
	 	 	 1777  : out <= -3420;
	 	 	 1778  : out <= -3418;
	 	 	 1779  : out <= -3415;
	 	 	 1780  : out <= -3413;
	 	 	 1781  : out <= -3411;
	 	 	 1782  : out <= -3408;
	 	 	 1783  : out <= -3406;
	 	 	 1784  : out <= -3404;
	 	 	 1785  : out <= -3402;
	 	 	 1786  : out <= -3399;
	 	 	 1787  : out <= -3397;
	 	 	 1788  : out <= -3395;
	 	 	 1789  : out <= -3392;
	 	 	 1790  : out <= -3390;
	 	 	 1791  : out <= -3388;
	 	 	 1792  : out <= -3386;
	 	 	 1793  : out <= -3383;
	 	 	 1794  : out <= -3381;
	 	 	 1795  : out <= -3379;
	 	 	 1796  : out <= -3376;
	 	 	 1797  : out <= -3374;
	 	 	 1798  : out <= -3372;
	 	 	 1799  : out <= -3370;
	 	 	 1800  : out <= -3367;
	 	 	 1801  : out <= -3365;
	 	 	 1802  : out <= -3363;
	 	 	 1803  : out <= -3361;
	 	 	 1804  : out <= -3358;
	 	 	 1805  : out <= -3356;
	 	 	 1806  : out <= -3354;
	 	 	 1807  : out <= -3351;
	 	 	 1808  : out <= -3349;
	 	 	 1809  : out <= -3347;
	 	 	 1810  : out <= -3345;
	 	 	 1811  : out <= -3342;
	 	 	 1812  : out <= -3340;
	 	 	 1813  : out <= -3338;
	 	 	 1814  : out <= -3336;
	 	 	 1815  : out <= -3333;
	 	 	 1816  : out <= -3331;
	 	 	 1817  : out <= -3329;
	 	 	 1818  : out <= -3327;
	 	 	 1819  : out <= -3324;
	 	 	 1820  : out <= -3322;
	 	 	 1821  : out <= -3320;
	 	 	 1822  : out <= -3318;
	 	 	 1823  : out <= -3315;
	 	 	 1824  : out <= -3313;
	 	 	 1825  : out <= -3311;
	 	 	 1826  : out <= -3309;
	 	 	 1827  : out <= -3306;
	 	 	 1828  : out <= -3304;
	 	 	 1829  : out <= -3302;
	 	 	 1830  : out <= -3300;
	 	 	 1831  : out <= -3297;
	 	 	 1832  : out <= -3295;
	 	 	 1833  : out <= -3293;
	 	 	 1834  : out <= -3291;
	 	 	 1835  : out <= -3288;
	 	 	 1836  : out <= -3286;
	 	 	 1837  : out <= -3284;
	 	 	 1838  : out <= -3282;
	 	 	 1839  : out <= -3280;
	 	 	 1840  : out <= -3277;
	 	 	 1841  : out <= -3275;
	 	 	 1842  : out <= -3273;
	 	 	 1843  : out <= -3271;
	 	 	 1844  : out <= -3268;
	 	 	 1845  : out <= -3266;
	 	 	 1846  : out <= -3264;
	 	 	 1847  : out <= -3262;
	 	 	 1848  : out <= -3260;
	 	 	 1849  : out <= -3257;
	 	 	 1850  : out <= -3255;
	 	 	 1851  : out <= -3253;
	 	 	 1852  : out <= -3251;
	 	 	 1853  : out <= -3248;
	 	 	 1854  : out <= -3246;
	 	 	 1855  : out <= -3244;
	 	 	 1856  : out <= -3242;
	 	 	 1857  : out <= -3240;
	 	 	 1858  : out <= -3237;
	 	 	 1859  : out <= -3235;
	 	 	 1860  : out <= -3233;
	 	 	 1861  : out <= -3231;
	 	 	 1862  : out <= -3229;
	 	 	 1863  : out <= -3226;
	 	 	 1864  : out <= -3224;
	 	 	 1865  : out <= -3222;
	 	 	 1866  : out <= -3220;
	 	 	 1867  : out <= -3218;
	 	 	 1868  : out <= -3215;
	 	 	 1869  : out <= -3213;
	 	 	 1870  : out <= -3211;
	 	 	 1871  : out <= -3209;
	 	 	 1872  : out <= -3207;
	 	 	 1873  : out <= -3204;
	 	 	 1874  : out <= -3202;
	 	 	 1875  : out <= -3200;
	 	 	 1876  : out <= -3198;
	 	 	 1877  : out <= -3196;
	 	 	 1878  : out <= -3194;
	 	 	 1879  : out <= -3191;
	 	 	 1880  : out <= -3189;
	 	 	 1881  : out <= -3187;
	 	 	 1882  : out <= -3185;
	 	 	 1883  : out <= -3183;
	 	 	 1884  : out <= -3181;
	 	 	 1885  : out <= -3178;
	 	 	 1886  : out <= -3176;
	 	 	 1887  : out <= -3174;
	 	 	 1888  : out <= -3172;
	 	 	 1889  : out <= -3170;
	 	 	 1890  : out <= -3167;
	 	 	 1891  : out <= -3165;
	 	 	 1892  : out <= -3163;
	 	 	 1893  : out <= -3161;
	 	 	 1894  : out <= -3159;
	 	 	 1895  : out <= -3157;
	 	 	 1896  : out <= -3155;
	 	 	 1897  : out <= -3152;
	 	 	 1898  : out <= -3150;
	 	 	 1899  : out <= -3148;
	 	 	 1900  : out <= -3146;
	 	 	 1901  : out <= -3144;
	 	 	 1902  : out <= -3142;
	 	 	 1903  : out <= -3139;
	 	 	 1904  : out <= -3137;
	 	 	 1905  : out <= -3135;
	 	 	 1906  : out <= -3133;
	 	 	 1907  : out <= -3131;
	 	 	 1908  : out <= -3129;
	 	 	 1909  : out <= -3127;
	 	 	 1910  : out <= -3124;
	 	 	 1911  : out <= -3122;
	 	 	 1912  : out <= -3120;
	 	 	 1913  : out <= -3118;
	 	 	 1914  : out <= -3116;
	 	 	 1915  : out <= -3114;
	 	 	 1916  : out <= -3112;
	 	 	 1917  : out <= -3109;
	 	 	 1918  : out <= -3107;
	 	 	 1919  : out <= -3105;
	 	 	 1920  : out <= -3103;
	 	 	 1921  : out <= -3101;
	 	 	 1922  : out <= -3099;
	 	 	 1923  : out <= -3097;
	 	 	 1924  : out <= -3094;
	 	 	 1925  : out <= -3092;
	 	 	 1926  : out <= -3090;
	 	 	 1927  : out <= -3088;
	 	 	 1928  : out <= -3086;
	 	 	 1929  : out <= -3084;
	 	 	 1930  : out <= -3082;
	 	 	 1931  : out <= -3080;
	 	 	 1932  : out <= -3077;
	 	 	 1933  : out <= -3075;
	 	 	 1934  : out <= -3073;
	 	 	 1935  : out <= -3071;
	 	 	 1936  : out <= -3069;
	 	 	 1937  : out <= -3067;
	 	 	 1938  : out <= -3065;
	 	 	 1939  : out <= -3063;
	 	 	 1940  : out <= -3061;
	 	 	 1941  : out <= -3058;
	 	 	 1942  : out <= -3056;
	 	 	 1943  : out <= -3054;
	 	 	 1944  : out <= -3052;
	 	 	 1945  : out <= -3050;
	 	 	 1946  : out <= -3048;
	 	 	 1947  : out <= -3046;
	 	 	 1948  : out <= -3044;
	 	 	 1949  : out <= -3042;
	 	 	 1950  : out <= -3039;
	 	 	 1951  : out <= -3037;
	 	 	 1952  : out <= -3035;
	 	 	 1953  : out <= -3033;
	 	 	 1954  : out <= -3031;
	 	 	 1955  : out <= -3029;
	 	 	 1956  : out <= -3027;
	 	 	 1957  : out <= -3025;
	 	 	 1958  : out <= -3023;
	 	 	 1959  : out <= -3021;
	 	 	 1960  : out <= -3019;
	 	 	 1961  : out <= -3016;
	 	 	 1962  : out <= -3014;
	 	 	 1963  : out <= -3012;
	 	 	 1964  : out <= -3010;
	 	 	 1965  : out <= -3008;
	 	 	 1966  : out <= -3006;
	 	 	 1967  : out <= -3004;
	 	 	 1968  : out <= -3002;
	 	 	 1969  : out <= -3000;
	 	 	 1970  : out <= -2998;
	 	 	 1971  : out <= -2996;
	 	 	 1972  : out <= -2994;
	 	 	 1973  : out <= -2991;
	 	 	 1974  : out <= -2989;
	 	 	 1975  : out <= -2987;
	 	 	 1976  : out <= -2985;
	 	 	 1977  : out <= -2983;
	 	 	 1978  : out <= -2981;
	 	 	 1979  : out <= -2979;
	 	 	 1980  : out <= -2977;
	 	 	 1981  : out <= -2975;
	 	 	 1982  : out <= -2973;
	 	 	 1983  : out <= -2971;
	 	 	 1984  : out <= -2969;
	 	 	 1985  : out <= -2967;
	 	 	 1986  : out <= -2965;
	 	 	 1987  : out <= -2962;
	 	 	 1988  : out <= -2960;
	 	 	 1989  : out <= -2958;
	 	 	 1990  : out <= -2956;
	 	 	 1991  : out <= -2954;
	 	 	 1992  : out <= -2952;
	 	 	 1993  : out <= -2950;
	 	 	 1994  : out <= -2948;
	 	 	 1995  : out <= -2946;
	 	 	 1996  : out <= -2944;
	 	 	 1997  : out <= -2942;
	 	 	 1998  : out <= -2940;
	 	 	 1999  : out <= -2938;
	 	 	 2000  : out <= -2936;
	 	 	 2001  : out <= -2934;
	 	 	 2002  : out <= -2932;
	 	 	 2003  : out <= -2930;
	 	 	 2004  : out <= -2928;
	 	 	 2005  : out <= -2926;
	 	 	 2006  : out <= -2924;
	 	 	 2007  : out <= -2921;
	 	 	 2008  : out <= -2919;
	 	 	 2009  : out <= -2917;
	 	 	 2010  : out <= -2915;
	 	 	 2011  : out <= -2913;
	 	 	 2012  : out <= -2911;
	 	 	 2013  : out <= -2909;
	 	 	 2014  : out <= -2907;
	 	 	 2015  : out <= -2905;
	 	 	 2016  : out <= -2903;
	 	 	 2017  : out <= -2901;
	 	 	 2018  : out <= -2899;
	 	 	 2019  : out <= -2897;
	 	 	 2020  : out <= -2895;
	 	 	 2021  : out <= -2893;
	 	 	 2022  : out <= -2891;
	 	 	 2023  : out <= -2889;
	 	 	 2024  : out <= -2887;
	 	 	 2025  : out <= -2885;
	 	 	 2026  : out <= -2883;
	 	 	 2027  : out <= -2881;
	 	 	 2028  : out <= -2879;
	 	 	 2029  : out <= -2877;
	 	 	 2030  : out <= -2875;
	 	 	 2031  : out <= -2873;
	 	 	 2032  : out <= -2871;
	 	 	 2033  : out <= -2869;
	 	 	 2034  : out <= -2867;
	 	 	 2035  : out <= -2865;
	 	 	 2036  : out <= -2863;
	 	 	 2037  : out <= -2861;
	 	 	 2038  : out <= -2859;
	 	 	 2039  : out <= -2857;
	 	 	 2040  : out <= -2855;
	 	 	 2041  : out <= -2853;
	 	 	 2042  : out <= -2851;
	 	 	 2043  : out <= -2849;
	 	 	 2044  : out <= -2847;
	 	 	 2045  : out <= -2845;
	 	 	 2046  : out <= -2843;
	 	 	 2047  : out <= -2841;
	 	 	 2048  : out <= -2839;
	 	 	 2049  : out <= -2837;
	 	 	 2050  : out <= -2835;
	 	 	 2051  : out <= -2833;
	 	 	 2052  : out <= -2831;
	 	 	 2053  : out <= -2829;
	 	 	 2054  : out <= -2827;
	 	 	 2055  : out <= -2825;
	 	 	 2056  : out <= -2823;
	 	 	 2057  : out <= -2821;
	 	 	 2058  : out <= -2819;
	 	 	 2059  : out <= -2817;
	 	 	 2060  : out <= -2815;
	 	 	 2061  : out <= -2813;
	 	 	 2062  : out <= -2811;
	 	 	 2063  : out <= -2809;
	 	 	 2064  : out <= -2807;
	 	 	 2065  : out <= -2805;
	 	 	 2066  : out <= -2803;
	 	 	 2067  : out <= -2801;
	 	 	 2068  : out <= -2799;
	 	 	 2069  : out <= -2797;
	 	 	 2070  : out <= -2795;
	 	 	 2071  : out <= -2793;
	 	 	 2072  : out <= -2791;
	 	 	 2073  : out <= -2789;
	 	 	 2074  : out <= -2787;
	 	 	 2075  : out <= -2785;
	 	 	 2076  : out <= -2783;
	 	 	 2077  : out <= -2781;
	 	 	 2078  : out <= -2779;
	 	 	 2079  : out <= -2777;
	 	 	 2080  : out <= -2775;
	 	 	 2081  : out <= -2773;
	 	 	 2082  : out <= -2771;
	 	 	 2083  : out <= -2769;
	 	 	 2084  : out <= -2767;
	 	 	 2085  : out <= -2765;
	 	 	 2086  : out <= -2763;
	 	 	 2087  : out <= -2761;
	 	 	 2088  : out <= -2759;
	 	 	 2089  : out <= -2757;
	 	 	 2090  : out <= -2755;
	 	 	 2091  : out <= -2754;
	 	 	 2092  : out <= -2752;
	 	 	 2093  : out <= -2750;
	 	 	 2094  : out <= -2748;
	 	 	 2095  : out <= -2746;
	 	 	 2096  : out <= -2744;
	 	 	 2097  : out <= -2742;
	 	 	 2098  : out <= -2740;
	 	 	 2099  : out <= -2738;
	 	 	 2100  : out <= -2736;
	 	 	 2101  : out <= -2734;
	 	 	 2102  : out <= -2732;
	 	 	 2103  : out <= -2730;
	 	 	 2104  : out <= -2728;
	 	 	 2105  : out <= -2726;
	 	 	 2106  : out <= -2724;
	 	 	 2107  : out <= -2722;
	 	 	 2108  : out <= -2720;
	 	 	 2109  : out <= -2718;
	 	 	 2110  : out <= -2716;
	 	 	 2111  : out <= -2715;
	 	 	 2112  : out <= -2713;
	 	 	 2113  : out <= -2711;
	 	 	 2114  : out <= -2709;
	 	 	 2115  : out <= -2707;
	 	 	 2116  : out <= -2705;
	 	 	 2117  : out <= -2703;
	 	 	 2118  : out <= -2701;
	 	 	 2119  : out <= -2699;
	 	 	 2120  : out <= -2697;
	 	 	 2121  : out <= -2695;
	 	 	 2122  : out <= -2693;
	 	 	 2123  : out <= -2691;
	 	 	 2124  : out <= -2689;
	 	 	 2125  : out <= -2687;
	 	 	 2126  : out <= -2686;
	 	 	 2127  : out <= -2684;
	 	 	 2128  : out <= -2682;
	 	 	 2129  : out <= -2680;
	 	 	 2130  : out <= -2678;
	 	 	 2131  : out <= -2676;
	 	 	 2132  : out <= -2674;
	 	 	 2133  : out <= -2672;
	 	 	 2134  : out <= -2670;
	 	 	 2135  : out <= -2668;
	 	 	 2136  : out <= -2666;
	 	 	 2137  : out <= -2664;
	 	 	 2138  : out <= -2662;
	 	 	 2139  : out <= -2661;
	 	 	 2140  : out <= -2659;
	 	 	 2141  : out <= -2657;
	 	 	 2142  : out <= -2655;
	 	 	 2143  : out <= -2653;
	 	 	 2144  : out <= -2651;
	 	 	 2145  : out <= -2649;
	 	 	 2146  : out <= -2647;
	 	 	 2147  : out <= -2645;
	 	 	 2148  : out <= -2643;
	 	 	 2149  : out <= -2641;
	 	 	 2150  : out <= -2640;
	 	 	 2151  : out <= -2638;
	 	 	 2152  : out <= -2636;
	 	 	 2153  : out <= -2634;
	 	 	 2154  : out <= -2632;
	 	 	 2155  : out <= -2630;
	 	 	 2156  : out <= -2628;
	 	 	 2157  : out <= -2626;
	 	 	 2158  : out <= -2624;
	 	 	 2159  : out <= -2622;
	 	 	 2160  : out <= -2621;
	 	 	 2161  : out <= -2619;
	 	 	 2162  : out <= -2617;
	 	 	 2163  : out <= -2615;
	 	 	 2164  : out <= -2613;
	 	 	 2165  : out <= -2611;
	 	 	 2166  : out <= -2609;
	 	 	 2167  : out <= -2607;
	 	 	 2168  : out <= -2605;
	 	 	 2169  : out <= -2604;
	 	 	 2170  : out <= -2602;
	 	 	 2171  : out <= -2600;
	 	 	 2172  : out <= -2598;
	 	 	 2173  : out <= -2596;
	 	 	 2174  : out <= -2594;
	 	 	 2175  : out <= -2592;
	 	 	 2176  : out <= -2590;
	 	 	 2177  : out <= -2588;
	 	 	 2178  : out <= -2587;
	 	 	 2179  : out <= -2585;
	 	 	 2180  : out <= -2583;
	 	 	 2181  : out <= -2581;
	 	 	 2182  : out <= -2579;
	 	 	 2183  : out <= -2577;
	 	 	 2184  : out <= -2575;
	 	 	 2185  : out <= -2573;
	 	 	 2186  : out <= -2572;
	 	 	 2187  : out <= -2570;
	 	 	 2188  : out <= -2568;
	 	 	 2189  : out <= -2566;
	 	 	 2190  : out <= -2564;
	 	 	 2191  : out <= -2562;
	 	 	 2192  : out <= -2560;
	 	 	 2193  : out <= -2558;
	 	 	 2194  : out <= -2557;
	 	 	 2195  : out <= -2555;
	 	 	 2196  : out <= -2553;
	 	 	 2197  : out <= -2551;
	 	 	 2198  : out <= -2549;
	 	 	 2199  : out <= -2547;
	 	 	 2200  : out <= -2545;
	 	 	 2201  : out <= -2544;
	 	 	 2202  : out <= -2542;
	 	 	 2203  : out <= -2540;
	 	 	 2204  : out <= -2538;
	 	 	 2205  : out <= -2536;
	 	 	 2206  : out <= -2534;
	 	 	 2207  : out <= -2532;
	 	 	 2208  : out <= -2531;
	 	 	 2209  : out <= -2529;
	 	 	 2210  : out <= -2527;
	 	 	 2211  : out <= -2525;
	 	 	 2212  : out <= -2523;
	 	 	 2213  : out <= -2521;
	 	 	 2214  : out <= -2519;
	 	 	 2215  : out <= -2518;
	 	 	 2216  : out <= -2516;
	 	 	 2217  : out <= -2514;
	 	 	 2218  : out <= -2512;
	 	 	 2219  : out <= -2510;
	 	 	 2220  : out <= -2508;
	 	 	 2221  : out <= -2506;
	 	 	 2222  : out <= -2505;
	 	 	 2223  : out <= -2503;
	 	 	 2224  : out <= -2501;
	 	 	 2225  : out <= -2499;
	 	 	 2226  : out <= -2497;
	 	 	 2227  : out <= -2495;
	 	 	 2228  : out <= -2494;
	 	 	 2229  : out <= -2492;
	 	 	 2230  : out <= -2490;
	 	 	 2231  : out <= -2488;
	 	 	 2232  : out <= -2486;
	 	 	 2233  : out <= -2484;
	 	 	 2234  : out <= -2483;
	 	 	 2235  : out <= -2481;
	 	 	 2236  : out <= -2479;
	 	 	 2237  : out <= -2477;
	 	 	 2238  : out <= -2475;
	 	 	 2239  : out <= -2473;
	 	 	 2240  : out <= -2472;
	 	 	 2241  : out <= -2470;
	 	 	 2242  : out <= -2468;
	 	 	 2243  : out <= -2466;
	 	 	 2244  : out <= -2464;
	 	 	 2245  : out <= -2462;
	 	 	 2246  : out <= -2461;
	 	 	 2247  : out <= -2459;
	 	 	 2248  : out <= -2457;
	 	 	 2249  : out <= -2455;
	 	 	 2250  : out <= -2453;
	 	 	 2251  : out <= -2452;
	 	 	 2252  : out <= -2450;
	 	 	 2253  : out <= -2448;
	 	 	 2254  : out <= -2446;
	 	 	 2255  : out <= -2444;
	 	 	 2256  : out <= -2442;
	 	 	 2257  : out <= -2441;
	 	 	 2258  : out <= -2439;
	 	 	 2259  : out <= -2437;
	 	 	 2260  : out <= -2435;
	 	 	 2261  : out <= -2433;
	 	 	 2262  : out <= -2432;
	 	 	 2263  : out <= -2430;
	 	 	 2264  : out <= -2428;
	 	 	 2265  : out <= -2426;
	 	 	 2266  : out <= -2424;
	 	 	 2267  : out <= -2423;
	 	 	 2268  : out <= -2421;
	 	 	 2269  : out <= -2419;
	 	 	 2270  : out <= -2417;
	 	 	 2271  : out <= -2415;
	 	 	 2272  : out <= -2413;
	 	 	 2273  : out <= -2412;
	 	 	 2274  : out <= -2410;
	 	 	 2275  : out <= -2408;
	 	 	 2276  : out <= -2406;
	 	 	 2277  : out <= -2404;
	 	 	 2278  : out <= -2403;
	 	 	 2279  : out <= -2401;
	 	 	 2280  : out <= -2399;
	 	 	 2281  : out <= -2397;
	 	 	 2282  : out <= -2395;
	 	 	 2283  : out <= -2394;
	 	 	 2284  : out <= -2392;
	 	 	 2285  : out <= -2390;
	 	 	 2286  : out <= -2388;
	 	 	 2287  : out <= -2387;
	 	 	 2288  : out <= -2385;
	 	 	 2289  : out <= -2383;
	 	 	 2290  : out <= -2381;
	 	 	 2291  : out <= -2379;
	 	 	 2292  : out <= -2378;
	 	 	 2293  : out <= -2376;
	 	 	 2294  : out <= -2374;
	 	 	 2295  : out <= -2372;
	 	 	 2296  : out <= -2370;
	 	 	 2297  : out <= -2369;
	 	 	 2298  : out <= -2367;
	 	 	 2299  : out <= -2365;
	 	 	 2300  : out <= -2363;
	 	 	 2301  : out <= -2362;
	 	 	 2302  : out <= -2360;
	 	 	 2303  : out <= -2358;
	 	 	 2304  : out <= -2356;
	 	 	 2305  : out <= -2354;
	 	 	 2306  : out <= -2353;
	 	 	 2307  : out <= -2351;
	 	 	 2308  : out <= -2349;
	 	 	 2309  : out <= -2347;
	 	 	 2310  : out <= -2346;
	 	 	 2311  : out <= -2344;
	 	 	 2312  : out <= -2342;
	 	 	 2313  : out <= -2340;
	 	 	 2314  : out <= -2338;
	 	 	 2315  : out <= -2337;
	 	 	 2316  : out <= -2335;
	 	 	 2317  : out <= -2333;
	 	 	 2318  : out <= -2331;
	 	 	 2319  : out <= -2330;
	 	 	 2320  : out <= -2328;
	 	 	 2321  : out <= -2326;
	 	 	 2322  : out <= -2324;
	 	 	 2323  : out <= -2323;
	 	 	 2324  : out <= -2321;
	 	 	 2325  : out <= -2319;
	 	 	 2326  : out <= -2317;
	 	 	 2327  : out <= -2316;
	 	 	 2328  : out <= -2314;
	 	 	 2329  : out <= -2312;
	 	 	 2330  : out <= -2310;
	 	 	 2331  : out <= -2308;
	 	 	 2332  : out <= -2307;
	 	 	 2333  : out <= -2305;
	 	 	 2334  : out <= -2303;
	 	 	 2335  : out <= -2301;
	 	 	 2336  : out <= -2300;
	 	 	 2337  : out <= -2298;
	 	 	 2338  : out <= -2296;
	 	 	 2339  : out <= -2294;
	 	 	 2340  : out <= -2293;
	 	 	 2341  : out <= -2291;
	 	 	 2342  : out <= -2289;
	 	 	 2343  : out <= -2287;
	 	 	 2344  : out <= -2286;
	 	 	 2345  : out <= -2284;
	 	 	 2346  : out <= -2282;
	 	 	 2347  : out <= -2280;
	 	 	 2348  : out <= -2279;
	 	 	 2349  : out <= -2277;
	 	 	 2350  : out <= -2275;
	 	 	 2351  : out <= -2273;
	 	 	 2352  : out <= -2272;
	 	 	 2353  : out <= -2270;
	 	 	 2354  : out <= -2268;
	 	 	 2355  : out <= -2267;
	 	 	 2356  : out <= -2265;
	 	 	 2357  : out <= -2263;
	 	 	 2358  : out <= -2261;
	 	 	 2359  : out <= -2260;
	 	 	 2360  : out <= -2258;
	 	 	 2361  : out <= -2256;
	 	 	 2362  : out <= -2254;
	 	 	 2363  : out <= -2253;
	 	 	 2364  : out <= -2251;
	 	 	 2365  : out <= -2249;
	 	 	 2366  : out <= -2247;
	 	 	 2367  : out <= -2246;
	 	 	 2368  : out <= -2244;
	 	 	 2369  : out <= -2242;
	 	 	 2370  : out <= -2241;
	 	 	 2371  : out <= -2239;
	 	 	 2372  : out <= -2237;
	 	 	 2373  : out <= -2235;
	 	 	 2374  : out <= -2234;
	 	 	 2375  : out <= -2232;
	 	 	 2376  : out <= -2230;
	 	 	 2377  : out <= -2228;
	 	 	 2378  : out <= -2227;
	 	 	 2379  : out <= -2225;
	 	 	 2380  : out <= -2223;
	 	 	 2381  : out <= -2222;
	 	 	 2382  : out <= -2220;
	 	 	 2383  : out <= -2218;
	 	 	 2384  : out <= -2216;
	 	 	 2385  : out <= -2215;
	 	 	 2386  : out <= -2213;
	 	 	 2387  : out <= -2211;
	 	 	 2388  : out <= -2210;
	 	 	 2389  : out <= -2208;
	 	 	 2390  : out <= -2206;
	 	 	 2391  : out <= -2204;
	 	 	 2392  : out <= -2203;
	 	 	 2393  : out <= -2201;
	 	 	 2394  : out <= -2199;
	 	 	 2395  : out <= -2198;
	 	 	 2396  : out <= -2196;
	 	 	 2397  : out <= -2194;
	 	 	 2398  : out <= -2192;
	 	 	 2399  : out <= -2191;
	 	 	 2400  : out <= -2189;
	 	 	 2401  : out <= -2187;
	 	 	 2402  : out <= -2186;
	 	 	 2403  : out <= -2184;
	 	 	 2404  : out <= -2182;
	 	 	 2405  : out <= -2180;
	 	 	 2406  : out <= -2179;
	 	 	 2407  : out <= -2177;
	 	 	 2408  : out <= -2175;
	 	 	 2409  : out <= -2174;
	 	 	 2410  : out <= -2172;
	 	 	 2411  : out <= -2170;
	 	 	 2412  : out <= -2169;
	 	 	 2413  : out <= -2167;
	 	 	 2414  : out <= -2165;
	 	 	 2415  : out <= -2163;
	 	 	 2416  : out <= -2162;
	 	 	 2417  : out <= -2160;
	 	 	 2418  : out <= -2158;
	 	 	 2419  : out <= -2157;
	 	 	 2420  : out <= -2155;
	 	 	 2421  : out <= -2153;
	 	 	 2422  : out <= -2152;
	 	 	 2423  : out <= -2150;
	 	 	 2424  : out <= -2148;
	 	 	 2425  : out <= -2147;
	 	 	 2426  : out <= -2145;
	 	 	 2427  : out <= -2143;
	 	 	 2428  : out <= -2141;
	 	 	 2429  : out <= -2140;
	 	 	 2430  : out <= -2138;
	 	 	 2431  : out <= -2136;
	 	 	 2432  : out <= -2135;
	 	 	 2433  : out <= -2133;
	 	 	 2434  : out <= -2131;
	 	 	 2435  : out <= -2130;
	 	 	 2436  : out <= -2128;
	 	 	 2437  : out <= -2126;
	 	 	 2438  : out <= -2125;
	 	 	 2439  : out <= -2123;
	 	 	 2440  : out <= -2121;
	 	 	 2441  : out <= -2120;
	 	 	 2442  : out <= -2118;
	 	 	 2443  : out <= -2116;
	 	 	 2444  : out <= -2115;
	 	 	 2445  : out <= -2113;
	 	 	 2446  : out <= -2111;
	 	 	 2447  : out <= -2110;
	 	 	 2448  : out <= -2108;
	 	 	 2449  : out <= -2106;
	 	 	 2450  : out <= -2105;
	 	 	 2451  : out <= -2103;
	 	 	 2452  : out <= -2101;
	 	 	 2453  : out <= -2100;
	 	 	 2454  : out <= -2098;
	 	 	 2455  : out <= -2096;
	 	 	 2456  : out <= -2095;
	 	 	 2457  : out <= -2093;
	 	 	 2458  : out <= -2091;
	 	 	 2459  : out <= -2090;
	 	 	 2460  : out <= -2088;
	 	 	 2461  : out <= -2086;
	 	 	 2462  : out <= -2085;
	 	 	 2463  : out <= -2083;
	 	 	 2464  : out <= -2081;
	 	 	 2465  : out <= -2080;
	 	 	 2466  : out <= -2078;
	 	 	 2467  : out <= -2076;
	 	 	 2468  : out <= -2075;
	 	 	 2469  : out <= -2073;
	 	 	 2470  : out <= -2071;
	 	 	 2471  : out <= -2070;
	 	 	 2472  : out <= -2068;
	 	 	 2473  : out <= -2066;
	 	 	 2474  : out <= -2065;
	 	 	 2475  : out <= -2063;
	 	 	 2476  : out <= -2061;
	 	 	 2477  : out <= -2060;
	 	 	 2478  : out <= -2058;
	 	 	 2479  : out <= -2056;
	 	 	 2480  : out <= -2055;
	 	 	 2481  : out <= -2053;
	 	 	 2482  : out <= -2051;
	 	 	 2483  : out <= -2050;
	 	 	 2484  : out <= -2048;
	 	 	 2485  : out <= -2046;
	 	 	 2486  : out <= -2045;
	 	 	 2487  : out <= -2043;
	 	 	 2488  : out <= -2041;
	 	 	 2489  : out <= -2040;
	 	 	 2490  : out <= -2038;
	 	 	 2491  : out <= -2037;
	 	 	 2492  : out <= -2035;
	 	 	 2493  : out <= -2033;
	 	 	 2494  : out <= -2032;
	 	 	 2495  : out <= -2030;
	 	 	 2496  : out <= -2028;
	 	 	 2497  : out <= -2027;
	 	 	 2498  : out <= -2025;
	 	 	 2499  : out <= -2023;
	 	 	 2500  : out <= -2022;
	 	 	 2501  : out <= -2020;
	 	 	 2502  : out <= -2019;
	 	 	 2503  : out <= -2017;
	 	 	 2504  : out <= -2015;
	 	 	 2505  : out <= -2014;
	 	 	 2506  : out <= -2012;
	 	 	 2507  : out <= -2010;
	 	 	 2508  : out <= -2009;
	 	 	 2509  : out <= -2007;
	 	 	 2510  : out <= -2005;
	 	 	 2511  : out <= -2004;
	 	 	 2512  : out <= -2002;
	 	 	 2513  : out <= -2001;
	 	 	 2514  : out <= -1999;
	 	 	 2515  : out <= -1997;
	 	 	 2516  : out <= -1996;
	 	 	 2517  : out <= -1994;
	 	 	 2518  : out <= -1992;
	 	 	 2519  : out <= -1991;
	 	 	 2520  : out <= -1989;
	 	 	 2521  : out <= -1988;
	 	 	 2522  : out <= -1986;
	 	 	 2523  : out <= -1984;
	 	 	 2524  : out <= -1983;
	 	 	 2525  : out <= -1981;
	 	 	 2526  : out <= -1979;
	 	 	 2527  : out <= -1978;
	 	 	 2528  : out <= -1976;
	 	 	 2529  : out <= -1975;
	 	 	 2530  : out <= -1973;
	 	 	 2531  : out <= -1971;
	 	 	 2532  : out <= -1970;
	 	 	 2533  : out <= -1968;
	 	 	 2534  : out <= -1966;
	 	 	 2535  : out <= -1965;
	 	 	 2536  : out <= -1963;
	 	 	 2537  : out <= -1962;
	 	 	 2538  : out <= -1960;
	 	 	 2539  : out <= -1958;
	 	 	 2540  : out <= -1957;
	 	 	 2541  : out <= -1955;
	 	 	 2542  : out <= -1954;
	 	 	 2543  : out <= -1952;
	 	 	 2544  : out <= -1950;
	 	 	 2545  : out <= -1949;
	 	 	 2546  : out <= -1947;
	 	 	 2547  : out <= -1945;
	 	 	 2548  : out <= -1944;
	 	 	 2549  : out <= -1942;
	 	 	 2550  : out <= -1941;
	 	 	 2551  : out <= -1939;
	 	 	 2552  : out <= -1937;
	 	 	 2553  : out <= -1936;
	 	 	 2554  : out <= -1934;
	 	 	 2555  : out <= -1933;
	 	 	 2556  : out <= -1931;
	 	 	 2557  : out <= -1929;
	 	 	 2558  : out <= -1928;
	 	 	 2559  : out <= -1926;
	 	 	 2560  : out <= -1925;
	 	 	 2561  : out <= -1923;
	 	 	 2562  : out <= -1921;
	 	 	 2563  : out <= -1920;
	 	 	 2564  : out <= -1918;
	 	 	 2565  : out <= -1917;
	 	 	 2566  : out <= -1915;
	 	 	 2567  : out <= -1913;
	 	 	 2568  : out <= -1912;
	 	 	 2569  : out <= -1910;
	 	 	 2570  : out <= -1909;
	 	 	 2571  : out <= -1907;
	 	 	 2572  : out <= -1905;
	 	 	 2573  : out <= -1904;
	 	 	 2574  : out <= -1902;
	 	 	 2575  : out <= -1901;
	 	 	 2576  : out <= -1899;
	 	 	 2577  : out <= -1898;
	 	 	 2578  : out <= -1896;
	 	 	 2579  : out <= -1894;
	 	 	 2580  : out <= -1893;
	 	 	 2581  : out <= -1891;
	 	 	 2582  : out <= -1890;
	 	 	 2583  : out <= -1888;
	 	 	 2584  : out <= -1886;
	 	 	 2585  : out <= -1885;
	 	 	 2586  : out <= -1883;
	 	 	 2587  : out <= -1882;
	 	 	 2588  : out <= -1880;
	 	 	 2589  : out <= -1878;
	 	 	 2590  : out <= -1877;
	 	 	 2591  : out <= -1875;
	 	 	 2592  : out <= -1874;
	 	 	 2593  : out <= -1872;
	 	 	 2594  : out <= -1871;
	 	 	 2595  : out <= -1869;
	 	 	 2596  : out <= -1867;
	 	 	 2597  : out <= -1866;
	 	 	 2598  : out <= -1864;
	 	 	 2599  : out <= -1863;
	 	 	 2600  : out <= -1861;
	 	 	 2601  : out <= -1860;
	 	 	 2602  : out <= -1858;
	 	 	 2603  : out <= -1856;
	 	 	 2604  : out <= -1855;
	 	 	 2605  : out <= -1853;
	 	 	 2606  : out <= -1852;
	 	 	 2607  : out <= -1850;
	 	 	 2608  : out <= -1849;
	 	 	 2609  : out <= -1847;
	 	 	 2610  : out <= -1845;
	 	 	 2611  : out <= -1844;
	 	 	 2612  : out <= -1842;
	 	 	 2613  : out <= -1841;
	 	 	 2614  : out <= -1839;
	 	 	 2615  : out <= -1838;
	 	 	 2616  : out <= -1836;
	 	 	 2617  : out <= -1834;
	 	 	 2618  : out <= -1833;
	 	 	 2619  : out <= -1831;
	 	 	 2620  : out <= -1830;
	 	 	 2621  : out <= -1828;
	 	 	 2622  : out <= -1827;
	 	 	 2623  : out <= -1825;
	 	 	 2624  : out <= -1823;
	 	 	 2625  : out <= -1822;
	 	 	 2626  : out <= -1820;
	 	 	 2627  : out <= -1819;
	 	 	 2628  : out <= -1817;
	 	 	 2629  : out <= -1816;
	 	 	 2630  : out <= -1814;
	 	 	 2631  : out <= -1813;
	 	 	 2632  : out <= -1811;
	 	 	 2633  : out <= -1809;
	 	 	 2634  : out <= -1808;
	 	 	 2635  : out <= -1806;
	 	 	 2636  : out <= -1805;
	 	 	 2637  : out <= -1803;
	 	 	 2638  : out <= -1802;
	 	 	 2639  : out <= -1800;
	 	 	 2640  : out <= -1799;
	 	 	 2641  : out <= -1797;
	 	 	 2642  : out <= -1795;
	 	 	 2643  : out <= -1794;
	 	 	 2644  : out <= -1792;
	 	 	 2645  : out <= -1791;
	 	 	 2646  : out <= -1789;
	 	 	 2647  : out <= -1788;
	 	 	 2648  : out <= -1786;
	 	 	 2649  : out <= -1785;
	 	 	 2650  : out <= -1783;
	 	 	 2651  : out <= -1782;
	 	 	 2652  : out <= -1780;
	 	 	 2653  : out <= -1778;
	 	 	 2654  : out <= -1777;
	 	 	 2655  : out <= -1775;
	 	 	 2656  : out <= -1774;
	 	 	 2657  : out <= -1772;
	 	 	 2658  : out <= -1771;
	 	 	 2659  : out <= -1769;
	 	 	 2660  : out <= -1768;
	 	 	 2661  : out <= -1766;
	 	 	 2662  : out <= -1765;
	 	 	 2663  : out <= -1763;
	 	 	 2664  : out <= -1762;
	 	 	 2665  : out <= -1760;
	 	 	 2666  : out <= -1758;
	 	 	 2667  : out <= -1757;
	 	 	 2668  : out <= -1755;
	 	 	 2669  : out <= -1754;
	 	 	 2670  : out <= -1752;
	 	 	 2671  : out <= -1751;
	 	 	 2672  : out <= -1749;
	 	 	 2673  : out <= -1748;
	 	 	 2674  : out <= -1746;
	 	 	 2675  : out <= -1745;
	 	 	 2676  : out <= -1743;
	 	 	 2677  : out <= -1742;
	 	 	 2678  : out <= -1740;
	 	 	 2679  : out <= -1739;
	 	 	 2680  : out <= -1737;
	 	 	 2681  : out <= -1735;
	 	 	 2682  : out <= -1734;
	 	 	 2683  : out <= -1732;
	 	 	 2684  : out <= -1731;
	 	 	 2685  : out <= -1729;
	 	 	 2686  : out <= -1728;
	 	 	 2687  : out <= -1726;
	 	 	 2688  : out <= -1725;
	 	 	 2689  : out <= -1723;
	 	 	 2690  : out <= -1722;
	 	 	 2691  : out <= -1720;
	 	 	 2692  : out <= -1719;
	 	 	 2693  : out <= -1717;
	 	 	 2694  : out <= -1716;
	 	 	 2695  : out <= -1714;
	 	 	 2696  : out <= -1713;
	 	 	 2697  : out <= -1711;
	 	 	 2698  : out <= -1710;
	 	 	 2699  : out <= -1708;
	 	 	 2700  : out <= -1707;
	 	 	 2701  : out <= -1705;
	 	 	 2702  : out <= -1704;
	 	 	 2703  : out <= -1702;
	 	 	 2704  : out <= -1700;
	 	 	 2705  : out <= -1699;
	 	 	 2706  : out <= -1697;
	 	 	 2707  : out <= -1696;
	 	 	 2708  : out <= -1694;
	 	 	 2709  : out <= -1693;
	 	 	 2710  : out <= -1691;
	 	 	 2711  : out <= -1690;
	 	 	 2712  : out <= -1688;
	 	 	 2713  : out <= -1687;
	 	 	 2714  : out <= -1685;
	 	 	 2715  : out <= -1684;
	 	 	 2716  : out <= -1682;
	 	 	 2717  : out <= -1681;
	 	 	 2718  : out <= -1679;
	 	 	 2719  : out <= -1678;
	 	 	 2720  : out <= -1676;
	 	 	 2721  : out <= -1675;
	 	 	 2722  : out <= -1673;
	 	 	 2723  : out <= -1672;
	 	 	 2724  : out <= -1670;
	 	 	 2725  : out <= -1669;
	 	 	 2726  : out <= -1667;
	 	 	 2727  : out <= -1666;
	 	 	 2728  : out <= -1664;
	 	 	 2729  : out <= -1663;
	 	 	 2730  : out <= -1661;
	 	 	 2731  : out <= -1660;
	 	 	 2732  : out <= -1658;
	 	 	 2733  : out <= -1657;
	 	 	 2734  : out <= -1655;
	 	 	 2735  : out <= -1654;
	 	 	 2736  : out <= -1652;
	 	 	 2737  : out <= -1651;
	 	 	 2738  : out <= -1649;
	 	 	 2739  : out <= -1648;
	 	 	 2740  : out <= -1646;
	 	 	 2741  : out <= -1645;
	 	 	 2742  : out <= -1643;
	 	 	 2743  : out <= -1642;
	 	 	 2744  : out <= -1640;
	 	 	 2745  : out <= -1639;
	 	 	 2746  : out <= -1637;
	 	 	 2747  : out <= -1636;
	 	 	 2748  : out <= -1634;
	 	 	 2749  : out <= -1633;
	 	 	 2750  : out <= -1631;
	 	 	 2751  : out <= -1630;
	 	 	 2752  : out <= -1628;
	 	 	 2753  : out <= -1627;
	 	 	 2754  : out <= -1625;
	 	 	 2755  : out <= -1624;
	 	 	 2756  : out <= -1622;
	 	 	 2757  : out <= -1621;
	 	 	 2758  : out <= -1619;
	 	 	 2759  : out <= -1618;
	 	 	 2760  : out <= -1617;
	 	 	 2761  : out <= -1615;
	 	 	 2762  : out <= -1614;
	 	 	 2763  : out <= -1612;
	 	 	 2764  : out <= -1611;
	 	 	 2765  : out <= -1609;
	 	 	 2766  : out <= -1608;
	 	 	 2767  : out <= -1606;
	 	 	 2768  : out <= -1605;
	 	 	 2769  : out <= -1603;
	 	 	 2770  : out <= -1602;
	 	 	 2771  : out <= -1600;
	 	 	 2772  : out <= -1599;
	 	 	 2773  : out <= -1597;
	 	 	 2774  : out <= -1596;
	 	 	 2775  : out <= -1594;
	 	 	 2776  : out <= -1593;
	 	 	 2777  : out <= -1591;
	 	 	 2778  : out <= -1590;
	 	 	 2779  : out <= -1588;
	 	 	 2780  : out <= -1587;
	 	 	 2781  : out <= -1585;
	 	 	 2782  : out <= -1584;
	 	 	 2783  : out <= -1583;
	 	 	 2784  : out <= -1581;
	 	 	 2785  : out <= -1580;
	 	 	 2786  : out <= -1578;
	 	 	 2787  : out <= -1577;
	 	 	 2788  : out <= -1575;
	 	 	 2789  : out <= -1574;
	 	 	 2790  : out <= -1572;
	 	 	 2791  : out <= -1571;
	 	 	 2792  : out <= -1569;
	 	 	 2793  : out <= -1568;
	 	 	 2794  : out <= -1566;
	 	 	 2795  : out <= -1565;
	 	 	 2796  : out <= -1563;
	 	 	 2797  : out <= -1562;
	 	 	 2798  : out <= -1561;
	 	 	 2799  : out <= -1559;
	 	 	 2800  : out <= -1558;
	 	 	 2801  : out <= -1556;
	 	 	 2802  : out <= -1555;
	 	 	 2803  : out <= -1553;
	 	 	 2804  : out <= -1552;
	 	 	 2805  : out <= -1550;
	 	 	 2806  : out <= -1549;
	 	 	 2807  : out <= -1547;
	 	 	 2808  : out <= -1546;
	 	 	 2809  : out <= -1544;
	 	 	 2810  : out <= -1543;
	 	 	 2811  : out <= -1542;
	 	 	 2812  : out <= -1540;
	 	 	 2813  : out <= -1539;
	 	 	 2814  : out <= -1537;
	 	 	 2815  : out <= -1536;
	 	 	 2816  : out <= -1534;
	 	 	 2817  : out <= -1533;
	 	 	 2818  : out <= -1531;
	 	 	 2819  : out <= -1530;
	 	 	 2820  : out <= -1528;
	 	 	 2821  : out <= -1527;
	 	 	 2822  : out <= -1526;
	 	 	 2823  : out <= -1524;
	 	 	 2824  : out <= -1523;
	 	 	 2825  : out <= -1521;
	 	 	 2826  : out <= -1520;
	 	 	 2827  : out <= -1518;
	 	 	 2828  : out <= -1517;
	 	 	 2829  : out <= -1515;
	 	 	 2830  : out <= -1514;
	 	 	 2831  : out <= -1512;
	 	 	 2832  : out <= -1511;
	 	 	 2833  : out <= -1510;
	 	 	 2834  : out <= -1508;
	 	 	 2835  : out <= -1507;
	 	 	 2836  : out <= -1505;
	 	 	 2837  : out <= -1504;
	 	 	 2838  : out <= -1502;
	 	 	 2839  : out <= -1501;
	 	 	 2840  : out <= -1499;
	 	 	 2841  : out <= -1498;
	 	 	 2842  : out <= -1497;
	 	 	 2843  : out <= -1495;
	 	 	 2844  : out <= -1494;
	 	 	 2845  : out <= -1492;
	 	 	 2846  : out <= -1491;
	 	 	 2847  : out <= -1489;
	 	 	 2848  : out <= -1488;
	 	 	 2849  : out <= -1487;
	 	 	 2850  : out <= -1485;
	 	 	 2851  : out <= -1484;
	 	 	 2852  : out <= -1482;
	 	 	 2853  : out <= -1481;
	 	 	 2854  : out <= -1479;
	 	 	 2855  : out <= -1478;
	 	 	 2856  : out <= -1476;
	 	 	 2857  : out <= -1475;
	 	 	 2858  : out <= -1474;
	 	 	 2859  : out <= -1472;
	 	 	 2860  : out <= -1471;
	 	 	 2861  : out <= -1469;
	 	 	 2862  : out <= -1468;
	 	 	 2863  : out <= -1466;
	 	 	 2864  : out <= -1465;
	 	 	 2865  : out <= -1464;
	 	 	 2866  : out <= -1462;
	 	 	 2867  : out <= -1461;
	 	 	 2868  : out <= -1459;
	 	 	 2869  : out <= -1458;
	 	 	 2870  : out <= -1456;
	 	 	 2871  : out <= -1455;
	 	 	 2872  : out <= -1454;
	 	 	 2873  : out <= -1452;
	 	 	 2874  : out <= -1451;
	 	 	 2875  : out <= -1449;
	 	 	 2876  : out <= -1448;
	 	 	 2877  : out <= -1446;
	 	 	 2878  : out <= -1445;
	 	 	 2879  : out <= -1444;
	 	 	 2880  : out <= -1442;
	 	 	 2881  : out <= -1441;
	 	 	 2882  : out <= -1439;
	 	 	 2883  : out <= -1438;
	 	 	 2884  : out <= -1437;
	 	 	 2885  : out <= -1435;
	 	 	 2886  : out <= -1434;
	 	 	 2887  : out <= -1432;
	 	 	 2888  : out <= -1431;
	 	 	 2889  : out <= -1429;
	 	 	 2890  : out <= -1428;
	 	 	 2891  : out <= -1427;
	 	 	 2892  : out <= -1425;
	 	 	 2893  : out <= -1424;
	 	 	 2894  : out <= -1422;
	 	 	 2895  : out <= -1421;
	 	 	 2896  : out <= -1420;
	 	 	 2897  : out <= -1418;
	 	 	 2898  : out <= -1417;
	 	 	 2899  : out <= -1415;
	 	 	 2900  : out <= -1414;
	 	 	 2901  : out <= -1412;
	 	 	 2902  : out <= -1411;
	 	 	 2903  : out <= -1410;
	 	 	 2904  : out <= -1408;
	 	 	 2905  : out <= -1407;
	 	 	 2906  : out <= -1405;
	 	 	 2907  : out <= -1404;
	 	 	 2908  : out <= -1403;
	 	 	 2909  : out <= -1401;
	 	 	 2910  : out <= -1400;
	 	 	 2911  : out <= -1398;
	 	 	 2912  : out <= -1397;
	 	 	 2913  : out <= -1396;
	 	 	 2914  : out <= -1394;
	 	 	 2915  : out <= -1393;
	 	 	 2916  : out <= -1391;
	 	 	 2917  : out <= -1390;
	 	 	 2918  : out <= -1389;
	 	 	 2919  : out <= -1387;
	 	 	 2920  : out <= -1386;
	 	 	 2921  : out <= -1384;
	 	 	 2922  : out <= -1383;
	 	 	 2923  : out <= -1381;
	 	 	 2924  : out <= -1380;
	 	 	 2925  : out <= -1379;
	 	 	 2926  : out <= -1377;
	 	 	 2927  : out <= -1376;
	 	 	 2928  : out <= -1374;
	 	 	 2929  : out <= -1373;
	 	 	 2930  : out <= -1372;
	 	 	 2931  : out <= -1370;
	 	 	 2932  : out <= -1369;
	 	 	 2933  : out <= -1368;
	 	 	 2934  : out <= -1366;
	 	 	 2935  : out <= -1365;
	 	 	 2936  : out <= -1363;
	 	 	 2937  : out <= -1362;
	 	 	 2938  : out <= -1361;
	 	 	 2939  : out <= -1359;
	 	 	 2940  : out <= -1358;
	 	 	 2941  : out <= -1356;
	 	 	 2942  : out <= -1355;
	 	 	 2943  : out <= -1354;
	 	 	 2944  : out <= -1352;
	 	 	 2945  : out <= -1351;
	 	 	 2946  : out <= -1349;
	 	 	 2947  : out <= -1348;
	 	 	 2948  : out <= -1347;
	 	 	 2949  : out <= -1345;
	 	 	 2950  : out <= -1344;
	 	 	 2951  : out <= -1342;
	 	 	 2952  : out <= -1341;
	 	 	 2953  : out <= -1340;
	 	 	 2954  : out <= -1338;
	 	 	 2955  : out <= -1337;
	 	 	 2956  : out <= -1336;
	 	 	 2957  : out <= -1334;
	 	 	 2958  : out <= -1333;
	 	 	 2959  : out <= -1331;
	 	 	 2960  : out <= -1330;
	 	 	 2961  : out <= -1329;
	 	 	 2962  : out <= -1327;
	 	 	 2963  : out <= -1326;
	 	 	 2964  : out <= -1324;
	 	 	 2965  : out <= -1323;
	 	 	 2966  : out <= -1322;
	 	 	 2967  : out <= -1320;
	 	 	 2968  : out <= -1319;
	 	 	 2969  : out <= -1318;
	 	 	 2970  : out <= -1316;
	 	 	 2971  : out <= -1315;
	 	 	 2972  : out <= -1313;
	 	 	 2973  : out <= -1312;
	 	 	 2974  : out <= -1311;
	 	 	 2975  : out <= -1309;
	 	 	 2976  : out <= -1308;
	 	 	 2977  : out <= -1307;
	 	 	 2978  : out <= -1305;
	 	 	 2979  : out <= -1304;
	 	 	 2980  : out <= -1302;
	 	 	 2981  : out <= -1301;
	 	 	 2982  : out <= -1300;
	 	 	 2983  : out <= -1298;
	 	 	 2984  : out <= -1297;
	 	 	 2985  : out <= -1296;
	 	 	 2986  : out <= -1294;
	 	 	 2987  : out <= -1293;
	 	 	 2988  : out <= -1291;
	 	 	 2989  : out <= -1290;
	 	 	 2990  : out <= -1289;
	 	 	 2991  : out <= -1287;
	 	 	 2992  : out <= -1286;
	 	 	 2993  : out <= -1285;
	 	 	 2994  : out <= -1283;
	 	 	 2995  : out <= -1282;
	 	 	 2996  : out <= -1280;
	 	 	 2997  : out <= -1279;
	 	 	 2998  : out <= -1278;
	 	 	 2999  : out <= -1276;
	 	 	 3000  : out <= -1275;
	 	 	 3001  : out <= -1274;
	 	 	 3002  : out <= -1272;
	 	 	 3003  : out <= -1271;
	 	 	 3004  : out <= -1270;
	 	 	 3005  : out <= -1268;
	 	 	 3006  : out <= -1267;
	 	 	 3007  : out <= -1265;
	 	 	 3008  : out <= -1264;
	 	 	 3009  : out <= -1263;
	 	 	 3010  : out <= -1261;
	 	 	 3011  : out <= -1260;
	 	 	 3012  : out <= -1259;
	 	 	 3013  : out <= -1257;
	 	 	 3014  : out <= -1256;
	 	 	 3015  : out <= -1255;
	 	 	 3016  : out <= -1253;
	 	 	 3017  : out <= -1252;
	 	 	 3018  : out <= -1250;
	 	 	 3019  : out <= -1249;
	 	 	 3020  : out <= -1248;
	 	 	 3021  : out <= -1246;
	 	 	 3022  : out <= -1245;
	 	 	 3023  : out <= -1244;
	 	 	 3024  : out <= -1242;
	 	 	 3025  : out <= -1241;
	 	 	 3026  : out <= -1240;
	 	 	 3027  : out <= -1238;
	 	 	 3028  : out <= -1237;
	 	 	 3029  : out <= -1236;
	 	 	 3030  : out <= -1234;
	 	 	 3031  : out <= -1233;
	 	 	 3032  : out <= -1232;
	 	 	 3033  : out <= -1230;
	 	 	 3034  : out <= -1229;
	 	 	 3035  : out <= -1227;
	 	 	 3036  : out <= -1226;
	 	 	 3037  : out <= -1225;
	 	 	 3038  : out <= -1223;
	 	 	 3039  : out <= -1222;
	 	 	 3040  : out <= -1221;
	 	 	 3041  : out <= -1219;
	 	 	 3042  : out <= -1218;
	 	 	 3043  : out <= -1217;
	 	 	 3044  : out <= -1215;
	 	 	 3045  : out <= -1214;
	 	 	 3046  : out <= -1213;
	 	 	 3047  : out <= -1211;
	 	 	 3048  : out <= -1210;
	 	 	 3049  : out <= -1209;
	 	 	 3050  : out <= -1207;
	 	 	 3051  : out <= -1206;
	 	 	 3052  : out <= -1205;
	 	 	 3053  : out <= -1203;
	 	 	 3054  : out <= -1202;
	 	 	 3055  : out <= -1201;
	 	 	 3056  : out <= -1199;
	 	 	 3057  : out <= -1198;
	 	 	 3058  : out <= -1197;
	 	 	 3059  : out <= -1195;
	 	 	 3060  : out <= -1194;
	 	 	 3061  : out <= -1193;
	 	 	 3062  : out <= -1191;
	 	 	 3063  : out <= -1190;
	 	 	 3064  : out <= -1189;
	 	 	 3065  : out <= -1187;
	 	 	 3066  : out <= -1186;
	 	 	 3067  : out <= -1185;
	 	 	 3068  : out <= -1183;
	 	 	 3069  : out <= -1182;
	 	 	 3070  : out <= -1181;
	 	 	 3071  : out <= -1179;
	 	 	 3072  : out <= -1178;
	 	 	 3073  : out <= -1177;
	 	 	 3074  : out <= -1175;
	 	 	 3075  : out <= -1174;
	 	 	 3076  : out <= -1173;
	 	 	 3077  : out <= -1171;
	 	 	 3078  : out <= -1170;
	 	 	 3079  : out <= -1169;
	 	 	 3080  : out <= -1167;
	 	 	 3081  : out <= -1166;
	 	 	 3082  : out <= -1165;
	 	 	 3083  : out <= -1163;
	 	 	 3084  : out <= -1162;
	 	 	 3085  : out <= -1161;
	 	 	 3086  : out <= -1159;
	 	 	 3087  : out <= -1158;
	 	 	 3088  : out <= -1157;
	 	 	 3089  : out <= -1155;
	 	 	 3090  : out <= -1154;
	 	 	 3091  : out <= -1153;
	 	 	 3092  : out <= -1151;
	 	 	 3093  : out <= -1150;
	 	 	 3094  : out <= -1149;
	 	 	 3095  : out <= -1147;
	 	 	 3096  : out <= -1146;
	 	 	 3097  : out <= -1145;
	 	 	 3098  : out <= -1143;
	 	 	 3099  : out <= -1142;
	 	 	 3100  : out <= -1141;
	 	 	 3101  : out <= -1139;
	 	 	 3102  : out <= -1138;
	 	 	 3103  : out <= -1137;
	 	 	 3104  : out <= -1135;
	 	 	 3105  : out <= -1134;
	 	 	 3106  : out <= -1133;
	 	 	 3107  : out <= -1131;
	 	 	 3108  : out <= -1130;
	 	 	 3109  : out <= -1129;
	 	 	 3110  : out <= -1127;
	 	 	 3111  : out <= -1126;
	 	 	 3112  : out <= -1125;
	 	 	 3113  : out <= -1124;
	 	 	 3114  : out <= -1122;
	 	 	 3115  : out <= -1121;
	 	 	 3116  : out <= -1120;
	 	 	 3117  : out <= -1118;
	 	 	 3118  : out <= -1117;
	 	 	 3119  : out <= -1116;
	 	 	 3120  : out <= -1114;
	 	 	 3121  : out <= -1113;
	 	 	 3122  : out <= -1112;
	 	 	 3123  : out <= -1110;
	 	 	 3124  : out <= -1109;
	 	 	 3125  : out <= -1108;
	 	 	 3126  : out <= -1106;
	 	 	 3127  : out <= -1105;
	 	 	 3128  : out <= -1104;
	 	 	 3129  : out <= -1103;
	 	 	 3130  : out <= -1101;
	 	 	 3131  : out <= -1100;
	 	 	 3132  : out <= -1099;
	 	 	 3133  : out <= -1097;
	 	 	 3134  : out <= -1096;
	 	 	 3135  : out <= -1095;
	 	 	 3136  : out <= -1093;
	 	 	 3137  : out <= -1092;
	 	 	 3138  : out <= -1091;
	 	 	 3139  : out <= -1089;
	 	 	 3140  : out <= -1088;
	 	 	 3141  : out <= -1087;
	 	 	 3142  : out <= -1086;
	 	 	 3143  : out <= -1084;
	 	 	 3144  : out <= -1083;
	 	 	 3145  : out <= -1082;
	 	 	 3146  : out <= -1080;
	 	 	 3147  : out <= -1079;
	 	 	 3148  : out <= -1078;
	 	 	 3149  : out <= -1076;
	 	 	 3150  : out <= -1075;
	 	 	 3151  : out <= -1074;
	 	 	 3152  : out <= -1073;
	 	 	 3153  : out <= -1071;
	 	 	 3154  : out <= -1070;
	 	 	 3155  : out <= -1069;
	 	 	 3156  : out <= -1067;
	 	 	 3157  : out <= -1066;
	 	 	 3158  : out <= -1065;
	 	 	 3159  : out <= -1063;
	 	 	 3160  : out <= -1062;
	 	 	 3161  : out <= -1061;
	 	 	 3162  : out <= -1060;
	 	 	 3163  : out <= -1058;
	 	 	 3164  : out <= -1057;
	 	 	 3165  : out <= -1056;
	 	 	 3166  : out <= -1054;
	 	 	 3167  : out <= -1053;
	 	 	 3168  : out <= -1052;
	 	 	 3169  : out <= -1051;
	 	 	 3170  : out <= -1049;
	 	 	 3171  : out <= -1048;
	 	 	 3172  : out <= -1047;
	 	 	 3173  : out <= -1045;
	 	 	 3174  : out <= -1044;
	 	 	 3175  : out <= -1043;
	 	 	 3176  : out <= -1041;
	 	 	 3177  : out <= -1040;
	 	 	 3178  : out <= -1039;
	 	 	 3179  : out <= -1038;
	 	 	 3180  : out <= -1036;
	 	 	 3181  : out <= -1035;
	 	 	 3182  : out <= -1034;
	 	 	 3183  : out <= -1032;
	 	 	 3184  : out <= -1031;
	 	 	 3185  : out <= -1030;
	 	 	 3186  : out <= -1029;
	 	 	 3187  : out <= -1027;
	 	 	 3188  : out <= -1026;
	 	 	 3189  : out <= -1025;
	 	 	 3190  : out <= -1023;
	 	 	 3191  : out <= -1022;
	 	 	 3192  : out <= -1021;
	 	 	 3193  : out <= -1020;
	 	 	 3194  : out <= -1018;
	 	 	 3195  : out <= -1017;
	 	 	 3196  : out <= -1016;
	 	 	 3197  : out <= -1014;
	 	 	 3198  : out <= -1013;
	 	 	 3199  : out <= -1012;
	 	 	 3200  : out <= -1011;
	 	 	 3201  : out <= -1009;
	 	 	 3202  : out <= -1008;
	 	 	 3203  : out <= -1007;
	 	 	 3204  : out <= -1006;
	 	 	 3205  : out <= -1004;
	 	 	 3206  : out <= -1003;
	 	 	 3207  : out <= -1002;
	 	 	 3208  : out <= -1000;
	 	 	 3209  : out <= -999;
	 	 	 3210  : out <= -998;
	 	 	 3211  : out <= -997;
	 	 	 3212  : out <= -995;
	 	 	 3213  : out <= -994;
	 	 	 3214  : out <= -993;
	 	 	 3215  : out <= -991;
	 	 	 3216  : out <= -990;
	 	 	 3217  : out <= -989;
	 	 	 3218  : out <= -988;
	 	 	 3219  : out <= -986;
	 	 	 3220  : out <= -985;
	 	 	 3221  : out <= -984;
	 	 	 3222  : out <= -983;
	 	 	 3223  : out <= -981;
	 	 	 3224  : out <= -980;
	 	 	 3225  : out <= -979;
	 	 	 3226  : out <= -977;
	 	 	 3227  : out <= -976;
	 	 	 3228  : out <= -975;
	 	 	 3229  : out <= -974;
	 	 	 3230  : out <= -972;
	 	 	 3231  : out <= -971;
	 	 	 3232  : out <= -970;
	 	 	 3233  : out <= -969;
	 	 	 3234  : out <= -967;
	 	 	 3235  : out <= -966;
	 	 	 3236  : out <= -965;
	 	 	 3237  : out <= -964;
	 	 	 3238  : out <= -962;
	 	 	 3239  : out <= -961;
	 	 	 3240  : out <= -960;
	 	 	 3241  : out <= -958;
	 	 	 3242  : out <= -957;
	 	 	 3243  : out <= -956;
	 	 	 3244  : out <= -955;
	 	 	 3245  : out <= -953;
	 	 	 3246  : out <= -952;
	 	 	 3247  : out <= -951;
	 	 	 3248  : out <= -950;
	 	 	 3249  : out <= -948;
	 	 	 3250  : out <= -947;
	 	 	 3251  : out <= -946;
	 	 	 3252  : out <= -945;
	 	 	 3253  : out <= -943;
	 	 	 3254  : out <= -942;
	 	 	 3255  : out <= -941;
	 	 	 3256  : out <= -940;
	 	 	 3257  : out <= -938;
	 	 	 3258  : out <= -937;
	 	 	 3259  : out <= -936;
	 	 	 3260  : out <= -935;
	 	 	 3261  : out <= -933;
	 	 	 3262  : out <= -932;
	 	 	 3263  : out <= -931;
	 	 	 3264  : out <= -930;
	 	 	 3265  : out <= -928;
	 	 	 3266  : out <= -927;
	 	 	 3267  : out <= -926;
	 	 	 3268  : out <= -925;
	 	 	 3269  : out <= -923;
	 	 	 3270  : out <= -922;
	 	 	 3271  : out <= -921;
	 	 	 3272  : out <= -920;
	 	 	 3273  : out <= -918;
	 	 	 3274  : out <= -917;
	 	 	 3275  : out <= -916;
	 	 	 3276  : out <= -914;
	 	 	 3277  : out <= -913;
	 	 	 3278  : out <= -912;
	 	 	 3279  : out <= -911;
	 	 	 3280  : out <= -909;
	 	 	 3281  : out <= -908;
	 	 	 3282  : out <= -907;
	 	 	 3283  : out <= -906;
	 	 	 3284  : out <= -905;
	 	 	 3285  : out <= -903;
	 	 	 3286  : out <= -902;
	 	 	 3287  : out <= -901;
	 	 	 3288  : out <= -900;
	 	 	 3289  : out <= -898;
	 	 	 3290  : out <= -897;
	 	 	 3291  : out <= -896;
	 	 	 3292  : out <= -895;
	 	 	 3293  : out <= -893;
	 	 	 3294  : out <= -892;
	 	 	 3295  : out <= -891;
	 	 	 3296  : out <= -890;
	 	 	 3297  : out <= -888;
	 	 	 3298  : out <= -887;
	 	 	 3299  : out <= -886;
	 	 	 3300  : out <= -885;
	 	 	 3301  : out <= -883;
	 	 	 3302  : out <= -882;
	 	 	 3303  : out <= -881;
	 	 	 3304  : out <= -880;
	 	 	 3305  : out <= -878;
	 	 	 3306  : out <= -877;
	 	 	 3307  : out <= -876;
	 	 	 3308  : out <= -875;
	 	 	 3309  : out <= -873;
	 	 	 3310  : out <= -872;
	 	 	 3311  : out <= -871;
	 	 	 3312  : out <= -870;
	 	 	 3313  : out <= -868;
	 	 	 3314  : out <= -867;
	 	 	 3315  : out <= -866;
	 	 	 3316  : out <= -865;
	 	 	 3317  : out <= -864;
	 	 	 3318  : out <= -862;
	 	 	 3319  : out <= -861;
	 	 	 3320  : out <= -860;
	 	 	 3321  : out <= -859;
	 	 	 3322  : out <= -857;
	 	 	 3323  : out <= -856;
	 	 	 3324  : out <= -855;
	 	 	 3325  : out <= -854;
	 	 	 3326  : out <= -852;
	 	 	 3327  : out <= -851;
	 	 	 3328  : out <= -850;
	 	 	 3329  : out <= -849;
	 	 	 3330  : out <= -848;
	 	 	 3331  : out <= -846;
	 	 	 3332  : out <= -845;
	 	 	 3333  : out <= -844;
	 	 	 3334  : out <= -843;
	 	 	 3335  : out <= -841;
	 	 	 3336  : out <= -840;
	 	 	 3337  : out <= -839;
	 	 	 3338  : out <= -838;
	 	 	 3339  : out <= -836;
	 	 	 3340  : out <= -835;
	 	 	 3341  : out <= -834;
	 	 	 3342  : out <= -833;
	 	 	 3343  : out <= -832;
	 	 	 3344  : out <= -830;
	 	 	 3345  : out <= -829;
	 	 	 3346  : out <= -828;
	 	 	 3347  : out <= -827;
	 	 	 3348  : out <= -825;
	 	 	 3349  : out <= -824;
	 	 	 3350  : out <= -823;
	 	 	 3351  : out <= -822;
	 	 	 3352  : out <= -821;
	 	 	 3353  : out <= -819;
	 	 	 3354  : out <= -818;
	 	 	 3355  : out <= -817;
	 	 	 3356  : out <= -816;
	 	 	 3357  : out <= -814;
	 	 	 3358  : out <= -813;
	 	 	 3359  : out <= -812;
	 	 	 3360  : out <= -811;
	 	 	 3361  : out <= -810;
	 	 	 3362  : out <= -808;
	 	 	 3363  : out <= -807;
	 	 	 3364  : out <= -806;
	 	 	 3365  : out <= -805;
	 	 	 3366  : out <= -803;
	 	 	 3367  : out <= -802;
	 	 	 3368  : out <= -801;
	 	 	 3369  : out <= -800;
	 	 	 3370  : out <= -799;
	 	 	 3371  : out <= -797;
	 	 	 3372  : out <= -796;
	 	 	 3373  : out <= -795;
	 	 	 3374  : out <= -794;
	 	 	 3375  : out <= -793;
	 	 	 3376  : out <= -791;
	 	 	 3377  : out <= -790;
	 	 	 3378  : out <= -789;
	 	 	 3379  : out <= -788;
	 	 	 3380  : out <= -786;
	 	 	 3381  : out <= -785;
	 	 	 3382  : out <= -784;
	 	 	 3383  : out <= -783;
	 	 	 3384  : out <= -782;
	 	 	 3385  : out <= -780;
	 	 	 3386  : out <= -779;
	 	 	 3387  : out <= -778;
	 	 	 3388  : out <= -777;
	 	 	 3389  : out <= -776;
	 	 	 3390  : out <= -774;
	 	 	 3391  : out <= -773;
	 	 	 3392  : out <= -772;
	 	 	 3393  : out <= -771;
	 	 	 3394  : out <= -770;
	 	 	 3395  : out <= -768;
	 	 	 3396  : out <= -767;
	 	 	 3397  : out <= -766;
	 	 	 3398  : out <= -765;
	 	 	 3399  : out <= -764;
	 	 	 3400  : out <= -762;
	 	 	 3401  : out <= -761;
	 	 	 3402  : out <= -760;
	 	 	 3403  : out <= -759;
	 	 	 3404  : out <= -758;
	 	 	 3405  : out <= -756;
	 	 	 3406  : out <= -755;
	 	 	 3407  : out <= -754;
	 	 	 3408  : out <= -753;
	 	 	 3409  : out <= -751;
	 	 	 3410  : out <= -750;
	 	 	 3411  : out <= -749;
	 	 	 3412  : out <= -748;
	 	 	 3413  : out <= -747;
	 	 	 3414  : out <= -745;
	 	 	 3415  : out <= -744;
	 	 	 3416  : out <= -743;
	 	 	 3417  : out <= -742;
	 	 	 3418  : out <= -741;
	 	 	 3419  : out <= -739;
	 	 	 3420  : out <= -738;
	 	 	 3421  : out <= -737;
	 	 	 3422  : out <= -736;
	 	 	 3423  : out <= -735;
	 	 	 3424  : out <= -734;
	 	 	 3425  : out <= -732;
	 	 	 3426  : out <= -731;
	 	 	 3427  : out <= -730;
	 	 	 3428  : out <= -729;
	 	 	 3429  : out <= -728;
	 	 	 3430  : out <= -726;
	 	 	 3431  : out <= -725;
	 	 	 3432  : out <= -724;
	 	 	 3433  : out <= -723;
	 	 	 3434  : out <= -722;
	 	 	 3435  : out <= -720;
	 	 	 3436  : out <= -719;
	 	 	 3437  : out <= -718;
	 	 	 3438  : out <= -717;
	 	 	 3439  : out <= -716;
	 	 	 3440  : out <= -714;
	 	 	 3441  : out <= -713;
	 	 	 3442  : out <= -712;
	 	 	 3443  : out <= -711;
	 	 	 3444  : out <= -710;
	 	 	 3445  : out <= -708;
	 	 	 3446  : out <= -707;
	 	 	 3447  : out <= -706;
	 	 	 3448  : out <= -705;
	 	 	 3449  : out <= -704;
	 	 	 3450  : out <= -703;
	 	 	 3451  : out <= -701;
	 	 	 3452  : out <= -700;
	 	 	 3453  : out <= -699;
	 	 	 3454  : out <= -698;
	 	 	 3455  : out <= -697;
	 	 	 3456  : out <= -695;
	 	 	 3457  : out <= -694;
	 	 	 3458  : out <= -693;
	 	 	 3459  : out <= -692;
	 	 	 3460  : out <= -691;
	 	 	 3461  : out <= -689;
	 	 	 3462  : out <= -688;
	 	 	 3463  : out <= -687;
	 	 	 3464  : out <= -686;
	 	 	 3465  : out <= -685;
	 	 	 3466  : out <= -684;
	 	 	 3467  : out <= -682;
	 	 	 3468  : out <= -681;
	 	 	 3469  : out <= -680;
	 	 	 3470  : out <= -679;
	 	 	 3471  : out <= -678;
	 	 	 3472  : out <= -676;
	 	 	 3473  : out <= -675;
	 	 	 3474  : out <= -674;
	 	 	 3475  : out <= -673;
	 	 	 3476  : out <= -672;
	 	 	 3477  : out <= -671;
	 	 	 3478  : out <= -669;
	 	 	 3479  : out <= -668;
	 	 	 3480  : out <= -667;
	 	 	 3481  : out <= -666;
	 	 	 3482  : out <= -665;
	 	 	 3483  : out <= -664;
	 	 	 3484  : out <= -662;
	 	 	 3485  : out <= -661;
	 	 	 3486  : out <= -660;
	 	 	 3487  : out <= -659;
	 	 	 3488  : out <= -658;
	 	 	 3489  : out <= -656;
	 	 	 3490  : out <= -655;
	 	 	 3491  : out <= -654;
	 	 	 3492  : out <= -653;
	 	 	 3493  : out <= -652;
	 	 	 3494  : out <= -651;
	 	 	 3495  : out <= -649;
	 	 	 3496  : out <= -648;
	 	 	 3497  : out <= -647;
	 	 	 3498  : out <= -646;
	 	 	 3499  : out <= -645;
	 	 	 3500  : out <= -644;
	 	 	 3501  : out <= -642;
	 	 	 3502  : out <= -641;
	 	 	 3503  : out <= -640;
	 	 	 3504  : out <= -639;
	 	 	 3505  : out <= -638;
	 	 	 3506  : out <= -637;
	 	 	 3507  : out <= -635;
	 	 	 3508  : out <= -634;
	 	 	 3509  : out <= -633;
	 	 	 3510  : out <= -632;
	 	 	 3511  : out <= -631;
	 	 	 3512  : out <= -630;
	 	 	 3513  : out <= -628;
	 	 	 3514  : out <= -627;
	 	 	 3515  : out <= -626;
	 	 	 3516  : out <= -625;
	 	 	 3517  : out <= -624;
	 	 	 3518  : out <= -623;
	 	 	 3519  : out <= -621;
	 	 	 3520  : out <= -620;
	 	 	 3521  : out <= -619;
	 	 	 3522  : out <= -618;
	 	 	 3523  : out <= -617;
	 	 	 3524  : out <= -616;
	 	 	 3525  : out <= -614;
	 	 	 3526  : out <= -613;
	 	 	 3527  : out <= -612;
	 	 	 3528  : out <= -611;
	 	 	 3529  : out <= -610;
	 	 	 3530  : out <= -609;
	 	 	 3531  : out <= -607;
	 	 	 3532  : out <= -606;
	 	 	 3533  : out <= -605;
	 	 	 3534  : out <= -604;
	 	 	 3535  : out <= -603;
	 	 	 3536  : out <= -602;
	 	 	 3537  : out <= -601;
	 	 	 3538  : out <= -599;
	 	 	 3539  : out <= -598;
	 	 	 3540  : out <= -597;
	 	 	 3541  : out <= -596;
	 	 	 3542  : out <= -595;
	 	 	 3543  : out <= -594;
	 	 	 3544  : out <= -592;
	 	 	 3545  : out <= -591;
	 	 	 3546  : out <= -590;
	 	 	 3547  : out <= -589;
	 	 	 3548  : out <= -588;
	 	 	 3549  : out <= -587;
	 	 	 3550  : out <= -585;
	 	 	 3551  : out <= -584;
	 	 	 3552  : out <= -583;
	 	 	 3553  : out <= -582;
	 	 	 3554  : out <= -581;
	 	 	 3555  : out <= -580;
	 	 	 3556  : out <= -579;
	 	 	 3557  : out <= -577;
	 	 	 3558  : out <= -576;
	 	 	 3559  : out <= -575;
	 	 	 3560  : out <= -574;
	 	 	 3561  : out <= -573;
	 	 	 3562  : out <= -572;
	 	 	 3563  : out <= -571;
	 	 	 3564  : out <= -569;
	 	 	 3565  : out <= -568;
	 	 	 3566  : out <= -567;
	 	 	 3567  : out <= -566;
	 	 	 3568  : out <= -565;
	 	 	 3569  : out <= -564;
	 	 	 3570  : out <= -562;
	 	 	 3571  : out <= -561;
	 	 	 3572  : out <= -560;
	 	 	 3573  : out <= -559;
	 	 	 3574  : out <= -558;
	 	 	 3575  : out <= -557;
	 	 	 3576  : out <= -556;
	 	 	 3577  : out <= -554;
	 	 	 3578  : out <= -553;
	 	 	 3579  : out <= -552;
	 	 	 3580  : out <= -551;
	 	 	 3581  : out <= -550;
	 	 	 3582  : out <= -549;
	 	 	 3583  : out <= -548;
	 	 	 3584  : out <= -546;
	 	 	 3585  : out <= -545;
	 	 	 3586  : out <= -544;
	 	 	 3587  : out <= -543;
	 	 	 3588  : out <= -542;
	 	 	 3589  : out <= -541;
	 	 	 3590  : out <= -540;
	 	 	 3591  : out <= -538;
	 	 	 3592  : out <= -537;
	 	 	 3593  : out <= -536;
	 	 	 3594  : out <= -535;
	 	 	 3595  : out <= -534;
	 	 	 3596  : out <= -533;
	 	 	 3597  : out <= -532;
	 	 	 3598  : out <= -530;
	 	 	 3599  : out <= -529;
	 	 	 3600  : out <= -528;
	 	 	 3601  : out <= -527;
	 	 	 3602  : out <= -526;
	 	 	 3603  : out <= -525;
	 	 	 3604  : out <= -524;
	 	 	 3605  : out <= -523;
	 	 	 3606  : out <= -521;
	 	 	 3607  : out <= -520;
	 	 	 3608  : out <= -519;
	 	 	 3609  : out <= -518;
	 	 	 3610  : out <= -517;
	 	 	 3611  : out <= -516;
	 	 	 3612  : out <= -515;
	 	 	 3613  : out <= -513;
	 	 	 3614  : out <= -512;
	 	 	 3615  : out <= -511;
	 	 	 3616  : out <= -510;
	 	 	 3617  : out <= -509;
	 	 	 3618  : out <= -508;
	 	 	 3619  : out <= -507;
	 	 	 3620  : out <= -506;
	 	 	 3621  : out <= -504;
	 	 	 3622  : out <= -503;
	 	 	 3623  : out <= -502;
	 	 	 3624  : out <= -501;
	 	 	 3625  : out <= -500;
	 	 	 3626  : out <= -499;
	 	 	 3627  : out <= -498;
	 	 	 3628  : out <= -496;
	 	 	 3629  : out <= -495;
	 	 	 3630  : out <= -494;
	 	 	 3631  : out <= -493;
	 	 	 3632  : out <= -492;
	 	 	 3633  : out <= -491;
	 	 	 3634  : out <= -490;
	 	 	 3635  : out <= -489;
	 	 	 3636  : out <= -487;
	 	 	 3637  : out <= -486;
	 	 	 3638  : out <= -485;
	 	 	 3639  : out <= -484;
	 	 	 3640  : out <= -483;
	 	 	 3641  : out <= -482;
	 	 	 3642  : out <= -481;
	 	 	 3643  : out <= -480;
	 	 	 3644  : out <= -478;
	 	 	 3645  : out <= -477;
	 	 	 3646  : out <= -476;
	 	 	 3647  : out <= -475;
	 	 	 3648  : out <= -474;
	 	 	 3649  : out <= -473;
	 	 	 3650  : out <= -472;
	 	 	 3651  : out <= -471;
	 	 	 3652  : out <= -469;
	 	 	 3653  : out <= -468;
	 	 	 3654  : out <= -467;
	 	 	 3655  : out <= -466;
	 	 	 3656  : out <= -465;
	 	 	 3657  : out <= -464;
	 	 	 3658  : out <= -463;
	 	 	 3659  : out <= -462;
	 	 	 3660  : out <= -460;
	 	 	 3661  : out <= -459;
	 	 	 3662  : out <= -458;
	 	 	 3663  : out <= -457;
	 	 	 3664  : out <= -456;
	 	 	 3665  : out <= -455;
	 	 	 3666  : out <= -454;
	 	 	 3667  : out <= -453;
	 	 	 3668  : out <= -452;
	 	 	 3669  : out <= -450;
	 	 	 3670  : out <= -449;
	 	 	 3671  : out <= -448;
	 	 	 3672  : out <= -447;
	 	 	 3673  : out <= -446;
	 	 	 3674  : out <= -445;
	 	 	 3675  : out <= -444;
	 	 	 3676  : out <= -443;
	 	 	 3677  : out <= -442;
	 	 	 3678  : out <= -440;
	 	 	 3679  : out <= -439;
	 	 	 3680  : out <= -438;
	 	 	 3681  : out <= -437;
	 	 	 3682  : out <= -436;
	 	 	 3683  : out <= -435;
	 	 	 3684  : out <= -434;
	 	 	 3685  : out <= -433;
	 	 	 3686  : out <= -432;
	 	 	 3687  : out <= -430;
	 	 	 3688  : out <= -429;
	 	 	 3689  : out <= -428;
	 	 	 3690  : out <= -427;
	 	 	 3691  : out <= -426;
	 	 	 3692  : out <= -425;
	 	 	 3693  : out <= -424;
	 	 	 3694  : out <= -423;
	 	 	 3695  : out <= -422;
	 	 	 3696  : out <= -420;
	 	 	 3697  : out <= -419;
	 	 	 3698  : out <= -418;
	 	 	 3699  : out <= -417;
	 	 	 3700  : out <= -416;
	 	 	 3701  : out <= -415;
	 	 	 3702  : out <= -414;
	 	 	 3703  : out <= -413;
	 	 	 3704  : out <= -412;
	 	 	 3705  : out <= -410;
	 	 	 3706  : out <= -409;
	 	 	 3707  : out <= -408;
	 	 	 3708  : out <= -407;
	 	 	 3709  : out <= -406;
	 	 	 3710  : out <= -405;
	 	 	 3711  : out <= -404;
	 	 	 3712  : out <= -403;
	 	 	 3713  : out <= -402;
	 	 	 3714  : out <= -401;
	 	 	 3715  : out <= -399;
	 	 	 3716  : out <= -398;
	 	 	 3717  : out <= -397;
	 	 	 3718  : out <= -396;
	 	 	 3719  : out <= -395;
	 	 	 3720  : out <= -394;
	 	 	 3721  : out <= -393;
	 	 	 3722  : out <= -392;
	 	 	 3723  : out <= -391;
	 	 	 3724  : out <= -389;
	 	 	 3725  : out <= -388;
	 	 	 3726  : out <= -387;
	 	 	 3727  : out <= -386;
	 	 	 3728  : out <= -385;
	 	 	 3729  : out <= -384;
	 	 	 3730  : out <= -383;
	 	 	 3731  : out <= -382;
	 	 	 3732  : out <= -381;
	 	 	 3733  : out <= -380;
	 	 	 3734  : out <= -379;
	 	 	 3735  : out <= -377;
	 	 	 3736  : out <= -376;
	 	 	 3737  : out <= -375;
	 	 	 3738  : out <= -374;
	 	 	 3739  : out <= -373;
	 	 	 3740  : out <= -372;
	 	 	 3741  : out <= -371;
	 	 	 3742  : out <= -370;
	 	 	 3743  : out <= -369;
	 	 	 3744  : out <= -368;
	 	 	 3745  : out <= -366;
	 	 	 3746  : out <= -365;
	 	 	 3747  : out <= -364;
	 	 	 3748  : out <= -363;
	 	 	 3749  : out <= -362;
	 	 	 3750  : out <= -361;
	 	 	 3751  : out <= -360;
	 	 	 3752  : out <= -359;
	 	 	 3753  : out <= -358;
	 	 	 3754  : out <= -357;
	 	 	 3755  : out <= -356;
	 	 	 3756  : out <= -354;
	 	 	 3757  : out <= -353;
	 	 	 3758  : out <= -352;
	 	 	 3759  : out <= -351;
	 	 	 3760  : out <= -350;
	 	 	 3761  : out <= -349;
	 	 	 3762  : out <= -348;
	 	 	 3763  : out <= -347;
	 	 	 3764  : out <= -346;
	 	 	 3765  : out <= -345;
	 	 	 3766  : out <= -344;
	 	 	 3767  : out <= -342;
	 	 	 3768  : out <= -341;
	 	 	 3769  : out <= -340;
	 	 	 3770  : out <= -339;
	 	 	 3771  : out <= -338;
	 	 	 3772  : out <= -337;
	 	 	 3773  : out <= -336;
	 	 	 3774  : out <= -335;
	 	 	 3775  : out <= -334;
	 	 	 3776  : out <= -333;
	 	 	 3777  : out <= -332;
	 	 	 3778  : out <= -331;
	 	 	 3779  : out <= -329;
	 	 	 3780  : out <= -328;
	 	 	 3781  : out <= -327;
	 	 	 3782  : out <= -326;
	 	 	 3783  : out <= -325;
	 	 	 3784  : out <= -324;
	 	 	 3785  : out <= -323;
	 	 	 3786  : out <= -322;
	 	 	 3787  : out <= -321;
	 	 	 3788  : out <= -320;
	 	 	 3789  : out <= -319;
	 	 	 3790  : out <= -318;
	 	 	 3791  : out <= -316;
	 	 	 3792  : out <= -315;
	 	 	 3793  : out <= -314;
	 	 	 3794  : out <= -313;
	 	 	 3795  : out <= -312;
	 	 	 3796  : out <= -311;
	 	 	 3797  : out <= -310;
	 	 	 3798  : out <= -309;
	 	 	 3799  : out <= -308;
	 	 	 3800  : out <= -307;
	 	 	 3801  : out <= -306;
	 	 	 3802  : out <= -305;
	 	 	 3803  : out <= -304;
	 	 	 3804  : out <= -302;
	 	 	 3805  : out <= -301;
	 	 	 3806  : out <= -300;
	 	 	 3807  : out <= -299;
	 	 	 3808  : out <= -298;
	 	 	 3809  : out <= -297;
	 	 	 3810  : out <= -296;
	 	 	 3811  : out <= -295;
	 	 	 3812  : out <= -294;
	 	 	 3813  : out <= -293;
	 	 	 3814  : out <= -292;
	 	 	 3815  : out <= -291;
	 	 	 3816  : out <= -290;
	 	 	 3817  : out <= -288;
	 	 	 3818  : out <= -287;
	 	 	 3819  : out <= -286;
	 	 	 3820  : out <= -285;
	 	 	 3821  : out <= -284;
	 	 	 3822  : out <= -283;
	 	 	 3823  : out <= -282;
	 	 	 3824  : out <= -281;
	 	 	 3825  : out <= -280;
	 	 	 3826  : out <= -279;
	 	 	 3827  : out <= -278;
	 	 	 3828  : out <= -277;
	 	 	 3829  : out <= -276;
	 	 	 3830  : out <= -275;
	 	 	 3831  : out <= -273;
	 	 	 3832  : out <= -272;
	 	 	 3833  : out <= -271;
	 	 	 3834  : out <= -270;
	 	 	 3835  : out <= -269;
	 	 	 3836  : out <= -268;
	 	 	 3837  : out <= -267;
	 	 	 3838  : out <= -266;
	 	 	 3839  : out <= -265;
	 	 	 3840  : out <= -264;
	 	 	 3841  : out <= -263;
	 	 	 3842  : out <= -262;
	 	 	 3843  : out <= -261;
	 	 	 3844  : out <= -260;
	 	 	 3845  : out <= -259;
	 	 	 3846  : out <= -257;
	 	 	 3847  : out <= -256;
	 	 	 3848  : out <= -255;
	 	 	 3849  : out <= -254;
	 	 	 3850  : out <= -253;
	 	 	 3851  : out <= -252;
	 	 	 3852  : out <= -251;
	 	 	 3853  : out <= -250;
	 	 	 3854  : out <= -249;
	 	 	 3855  : out <= -248;
	 	 	 3856  : out <= -247;
	 	 	 3857  : out <= -246;
	 	 	 3858  : out <= -245;
	 	 	 3859  : out <= -244;
	 	 	 3860  : out <= -243;
	 	 	 3861  : out <= -242;
	 	 	 3862  : out <= -240;
	 	 	 3863  : out <= -239;
	 	 	 3864  : out <= -238;
	 	 	 3865  : out <= -237;
	 	 	 3866  : out <= -236;
	 	 	 3867  : out <= -235;
	 	 	 3868  : out <= -234;
	 	 	 3869  : out <= -233;
	 	 	 3870  : out <= -232;
	 	 	 3871  : out <= -231;
	 	 	 3872  : out <= -230;
	 	 	 3873  : out <= -229;
	 	 	 3874  : out <= -228;
	 	 	 3875  : out <= -227;
	 	 	 3876  : out <= -226;
	 	 	 3877  : out <= -225;
	 	 	 3878  : out <= -224;
	 	 	 3879  : out <= -222;
	 	 	 3880  : out <= -221;
	 	 	 3881  : out <= -220;
	 	 	 3882  : out <= -219;
	 	 	 3883  : out <= -218;
	 	 	 3884  : out <= -217;
	 	 	 3885  : out <= -216;
	 	 	 3886  : out <= -215;
	 	 	 3887  : out <= -214;
	 	 	 3888  : out <= -213;
	 	 	 3889  : out <= -212;
	 	 	 3890  : out <= -211;
	 	 	 3891  : out <= -210;
	 	 	 3892  : out <= -209;
	 	 	 3893  : out <= -208;
	 	 	 3894  : out <= -207;
	 	 	 3895  : out <= -206;
	 	 	 3896  : out <= -205;
	 	 	 3897  : out <= -203;
	 	 	 3898  : out <= -202;
	 	 	 3899  : out <= -201;
	 	 	 3900  : out <= -200;
	 	 	 3901  : out <= -199;
	 	 	 3902  : out <= -198;
	 	 	 3903  : out <= -197;
	 	 	 3904  : out <= -196;
	 	 	 3905  : out <= -195;
	 	 	 3906  : out <= -194;
	 	 	 3907  : out <= -193;
	 	 	 3908  : out <= -192;
	 	 	 3909  : out <= -191;
	 	 	 3910  : out <= -190;
	 	 	 3911  : out <= -189;
	 	 	 3912  : out <= -188;
	 	 	 3913  : out <= -187;
	 	 	 3914  : out <= -186;
	 	 	 3915  : out <= -185;
	 	 	 3916  : out <= -184;
	 	 	 3917  : out <= -183;
	 	 	 3918  : out <= -181;
	 	 	 3919  : out <= -180;
	 	 	 3920  : out <= -179;
	 	 	 3921  : out <= -178;
	 	 	 3922  : out <= -177;
	 	 	 3923  : out <= -176;
	 	 	 3924  : out <= -175;
	 	 	 3925  : out <= -174;
	 	 	 3926  : out <= -173;
	 	 	 3927  : out <= -172;
	 	 	 3928  : out <= -171;
	 	 	 3929  : out <= -170;
	 	 	 3930  : out <= -169;
	 	 	 3931  : out <= -168;
	 	 	 3932  : out <= -167;
	 	 	 3933  : out <= -166;
	 	 	 3934  : out <= -165;
	 	 	 3935  : out <= -164;
	 	 	 3936  : out <= -163;
	 	 	 3937  : out <= -162;
	 	 	 3938  : out <= -161;
	 	 	 3939  : out <= -160;
	 	 	 3940  : out <= -159;
	 	 	 3941  : out <= -158;
	 	 	 3942  : out <= -156;
	 	 	 3943  : out <= -155;
	 	 	 3944  : out <= -154;
	 	 	 3945  : out <= -153;
	 	 	 3946  : out <= -152;
	 	 	 3947  : out <= -151;
	 	 	 3948  : out <= -150;
	 	 	 3949  : out <= -149;
	 	 	 3950  : out <= -148;
	 	 	 3951  : out <= -147;
	 	 	 3952  : out <= -146;
	 	 	 3953  : out <= -145;
	 	 	 3954  : out <= -144;
	 	 	 3955  : out <= -143;
	 	 	 3956  : out <= -142;
	 	 	 3957  : out <= -141;
	 	 	 3958  : out <= -140;
	 	 	 3959  : out <= -139;
	 	 	 3960  : out <= -138;
	 	 	 3961  : out <= -137;
	 	 	 3962  : out <= -136;
	 	 	 3963  : out <= -135;
	 	 	 3964  : out <= -134;
	 	 	 3965  : out <= -133;
	 	 	 3966  : out <= -132;
	 	 	 3967  : out <= -131;
	 	 	 3968  : out <= -130;
	 	 	 3969  : out <= -129;
	 	 	 3970  : out <= -127;
	 	 	 3971  : out <= -126;
	 	 	 3972  : out <= -125;
	 	 	 3973  : out <= -124;
	 	 	 3974  : out <= -123;
	 	 	 3975  : out <= -122;
	 	 	 3976  : out <= -121;
	 	 	 3977  : out <= -120;
	 	 	 3978  : out <= -119;
	 	 	 3979  : out <= -118;
	 	 	 3980  : out <= -117;
	 	 	 3981  : out <= -116;
	 	 	 3982  : out <= -115;
	 	 	 3983  : out <= -114;
	 	 	 3984  : out <= -113;
	 	 	 3985  : out <= -112;
	 	 	 3986  : out <= -111;
	 	 	 3987  : out <= -110;
	 	 	 3988  : out <= -109;
	 	 	 3989  : out <= -108;
	 	 	 3990  : out <= -107;
	 	 	 3991  : out <= -106;
	 	 	 3992  : out <= -105;
	 	 	 3993  : out <= -104;
	 	 	 3994  : out <= -103;
	 	 	 3995  : out <= -102;
	 	 	 3996  : out <= -101;
	 	 	 3997  : out <= -100;
	 	 	 3998  : out <= -99;
	 	 	 3999  : out <= -98;
	 	 	 4000  : out <= -97;
	 	 	 4001  : out <= -96;
	 	 	 4002  : out <= -95;
	 	 	 4003  : out <= -94;
	 	 	 4004  : out <= -93;
	 	 	 4005  : out <= -92;
	 	 	 4006  : out <= -91;
	 	 	 4007  : out <= -89;
	 	 	 4008  : out <= -88;
	 	 	 4009  : out <= -87;
	 	 	 4010  : out <= -86;
	 	 	 4011  : out <= -85;
	 	 	 4012  : out <= -84;
	 	 	 4013  : out <= -83;
	 	 	 4014  : out <= -82;
	 	 	 4015  : out <= -81;
	 	 	 4016  : out <= -80;
	 	 	 4017  : out <= -79;
	 	 	 4018  : out <= -78;
	 	 	 4019  : out <= -77;
	 	 	 4020  : out <= -76;
	 	 	 4021  : out <= -75;
	 	 	 4022  : out <= -74;
	 	 	 4023  : out <= -73;
	 	 	 4024  : out <= -72;
	 	 	 4025  : out <= -71;
	 	 	 4026  : out <= -70;
	 	 	 4027  : out <= -69;
	 	 	 4028  : out <= -68;
	 	 	 4029  : out <= -67;
	 	 	 4030  : out <= -66;
	 	 	 4031  : out <= -65;
	 	 	 4032  : out <= -64;
	 	 	 4033  : out <= -63;
	 	 	 4034  : out <= -62;
	 	 	 4035  : out <= -61;
	 	 	 4036  : out <= -60;
	 	 	 4037  : out <= -59;
	 	 	 4038  : out <= -58;
	 	 	 4039  : out <= -57;
	 	 	 4040  : out <= -56;
	 	 	 4041  : out <= -55;
	 	 	 4042  : out <= -54;
	 	 	 4043  : out <= -53;
	 	 	 4044  : out <= -52;
	 	 	 4045  : out <= -51;
	 	 	 4046  : out <= -50;
	 	 	 4047  : out <= -49;
	 	 	 4048  : out <= -48;
	 	 	 4049  : out <= -47;
	 	 	 4050  : out <= -46;
	 	 	 4051  : out <= -45;
	 	 	 4052  : out <= -44;
	 	 	 4053  : out <= -43;
	 	 	 4054  : out <= -42;
	 	 	 4055  : out <= -41;
	 	 	 4056  : out <= -40;
	 	 	 4057  : out <= -39;
	 	 	 4058  : out <= -38;
	 	 	 4059  : out <= -37;
	 	 	 4060  : out <= -36;
	 	 	 4061  : out <= -35;
	 	 	 4062  : out <= -34;
	 	 	 4063  : out <= -33;
	 	 	 4064  : out <= -32;
	 	 	 4065  : out <= -31;
	 	 	 4066  : out <= -30;
	 	 	 4067  : out <= -29;
	 	 	 4068  : out <= -28;
	 	 	 4069  : out <= -27;
	 	 	 4070  : out <= -26;
	 	 	 4071  : out <= -25;
	 	 	 4072  : out <= -24;
	 	 	 4073  : out <= -23;
	 	 	 4074  : out <= -22;
	 	 	 4075  : out <= -21;
	 	 	 4076  : out <= -20;
	 	 	 4077  : out <= -19;
	 	 	 4078  : out <= -18;
	 	 	 4079  : out <= -17;
	 	 	 4080  : out <= -16;
	 	 	 4081  : out <= -15;
	 	 	 4082  : out <= -14;
	 	 	 4083  : out <= -13;
	 	 	 4084  : out <= -12;
	 	 	 4085  : out <= -11;
	 	 	 4086  : out <= -10;
	 	 	 4087  : out <= -9;
	 	 	 4088  : out <= -8;
	 	 	 4089  : out <= -7;
	 	 	 4090  : out <= -6;
	 	 	 4091  : out <= -5;
	 	 	 4092  : out <= -4;
	 	 	 4093  : out <= -3;
	 	 	 4094  : out <= -2;
	 	 	 4095  : out <= -1;
	 	 	 4096  : out <= 0;
	 	 	 default : out <= 0;
	 	 endcase
	 endmodule
