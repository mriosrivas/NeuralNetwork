//ROWS = output neurons
//COLUMNS = input size

// 3 -> 4 -> 2 -> 1


`ifndef forward_net_header
`define forward_net_header
    parameter L1 = 3; // Number of Rows
    parameter L2 = 4; // Number of Columns
    parameter L3 = 2;
    parameter L4 = 1;
`endif
