module sigma_int(input logic [15:0] in,
	 output logic [11:0] out);
	 	 always_comb
	 	 	 if (in >= 0 && in <= 2) out = 2047;
	 	 	 else if (in >= 3 && in <= 6) out = 2048;
	 	 	 else if (in >= 7 && in <= 10) out = 2049;
	 	 	 else if (in >= 11 && in <= 14) out = 2050;
	 	 	 else if (in >= 15 && in <= 18) out = 2051;
	 	 	 else if (in >= 19 && in <= 22) out = 2052;
	 	 	 else if (in >= 23 && in <= 26) out = 2053;
	 	 	 else if (in >= 27 && in <= 30) out = 2054;
	 	 	 else if (in >= 31 && in <= 34) out = 2055;
	 	 	 else if (in >= 35 && in <= 38) out = 2056;
	 	 	 else if (in >= 39 && in <= 42) out = 2057;
	 	 	 else if (in >= 43 && in <= 46) out = 2058;
	 	 	 else if (in >= 47 && in <= 50) out = 2059;
	 	 	 else if (in >= 51 && in <= 54) out = 2060;
	 	 	 else if (in >= 55 && in <= 58) out = 2061;
	 	 	 else if (in >= 59 && in <= 62) out = 2062;
	 	 	 else if (in >= 63 && in <= 66) out = 2063;
	 	 	 else if (in >= 67 && in <= 70) out = 2064;
	 	 	 else if (in >= 71 && in <= 74) out = 2065;
	 	 	 else if (in >= 75 && in <= 78) out = 2066;
	 	 	 else if (in >= 79 && in <= 82) out = 2067;
	 	 	 else if (in >= 83 && in <= 86) out = 2068;
	 	 	 else if (in >= 87 && in <= 90) out = 2069;
	 	 	 else if (in >= 91 && in <= 94) out = 2070;
	 	 	 else if (in >= 95 && in <= 98) out = 2071;
	 	 	 else if (in >= 99 && in <= 102) out = 2072;
	 	 	 else if (in >= 103 && in <= 106) out = 2073;
	 	 	 else if (in >= 107 && in <= 110) out = 2074;
	 	 	 else if (in >= 111 && in <= 114) out = 2075;
	 	 	 else if (in >= 115 && in <= 118) out = 2076;
	 	 	 else if (in >= 119 && in <= 122) out = 2077;
	 	 	 else if (in >= 123 && in <= 126) out = 2078;
	 	 	 else if (in >= 127 && in <= 130) out = 2079;
	 	 	 else if (in >= 131 && in <= 134) out = 2080;
	 	 	 else if (in >= 135 && in <= 138) out = 2081;
	 	 	 else if (in >= 139 && in <= 142) out = 2082;
	 	 	 else if (in >= 143 && in <= 146) out = 2083;
	 	 	 else if (in >= 147 && in <= 150) out = 2084;
	 	 	 else if (in >= 151 && in <= 154) out = 2085;
	 	 	 else if (in >= 155 && in <= 158) out = 2086;
	 	 	 else if (in >= 159 && in <= 162) out = 2087;
	 	 	 else if (in >= 163 && in <= 166) out = 2088;
	 	 	 else if (in >= 167 && in <= 170) out = 2089;
	 	 	 else if (in >= 171 && in <= 174) out = 2090;
	 	 	 else if (in >= 175 && in <= 178) out = 2091;
	 	 	 else if (in >= 179 && in <= 182) out = 2092;
	 	 	 else if (in >= 183 && in <= 186) out = 2093;
	 	 	 else if (in >= 187 && in <= 190) out = 2094;
	 	 	 else if (in >= 191 && in <= 194) out = 2095;
	 	 	 else if (in >= 195 && in <= 198) out = 2096;
	 	 	 else if (in >= 199 && in <= 202) out = 2097;
	 	 	 else if (in >= 203 && in <= 206) out = 2098;
	 	 	 else if (in >= 207 && in <= 210) out = 2099;
	 	 	 else if (in >= 211 && in <= 214) out = 2100;
	 	 	 else if (in >= 215 && in <= 218) out = 2101;
	 	 	 else if (in >= 219 && in <= 222) out = 2102;
	 	 	 else if (in >= 223 && in <= 226) out = 2103;
	 	 	 else if (in >= 227 && in <= 230) out = 2104;
	 	 	 else if (in >= 231 && in <= 234) out = 2105;
	 	 	 else if (in >= 235 && in <= 238) out = 2106;
	 	 	 else if (in >= 239 && in <= 242) out = 2107;
	 	 	 else if (in >= 243 && in <= 246) out = 2108;
	 	 	 else if (in >= 247 && in <= 250) out = 2109;
	 	 	 else if (in >= 251 && in <= 254) out = 2110;
	 	 	 else if (in >= 255 && in <= 258) out = 2111;
	 	 	 else if (in >= 259 && in <= 262) out = 2112;
	 	 	 else if (in >= 263 && in <= 266) out = 2113;
	 	 	 else if (in >= 267 && in <= 270) out = 2114;
	 	 	 else if (in >= 271 && in <= 274) out = 2115;
	 	 	 else if (in >= 275 && in <= 278) out = 2116;
	 	 	 else if (in >= 279 && in <= 282) out = 2117;
	 	 	 else if (in >= 283 && in <= 286) out = 2118;
	 	 	 else if (in >= 287 && in <= 290) out = 2119;
	 	 	 else if (in >= 291 && in <= 294) out = 2120;
	 	 	 else if (in >= 295 && in <= 298) out = 2121;
	 	 	 else if (in >= 299 && in <= 302) out = 2122;
	 	 	 else if (in >= 303 && in <= 306) out = 2123;
	 	 	 else if (in >= 307 && in <= 310) out = 2124;
	 	 	 else if (in >= 311 && in <= 314) out = 2125;
	 	 	 else if (in >= 315 && in <= 318) out = 2126;
	 	 	 else if (in >= 319 && in <= 322) out = 2127;
	 	 	 else if (in >= 323 && in <= 326) out = 2128;
	 	 	 else if (in >= 327 && in <= 330) out = 2129;
	 	 	 else if (in >= 331 && in <= 334) out = 2130;
	 	 	 else if (in >= 335 && in <= 338) out = 2131;
	 	 	 else if (in >= 339 && in <= 342) out = 2132;
	 	 	 else if (in >= 343 && in <= 346) out = 2133;
	 	 	 else if (in >= 347 && in <= 350) out = 2134;
	 	 	 else if (in >= 351 && in <= 354) out = 2135;
	 	 	 else if (in >= 355 && in <= 358) out = 2136;
	 	 	 else if (in >= 359 && in <= 362) out = 2137;
	 	 	 else if (in >= 363 && in <= 366) out = 2138;
	 	 	 else if (in >= 367 && in <= 370) out = 2139;
	 	 	 else if (in >= 371 && in <= 374) out = 2140;
	 	 	 else if (in >= 375 && in <= 378) out = 2141;
	 	 	 else if (in >= 379 && in <= 382) out = 2142;
	 	 	 else if (in >= 383 && in <= 386) out = 2143;
	 	 	 else if (in >= 387 && in <= 390) out = 2144;
	 	 	 else if (in >= 391 && in <= 394) out = 2145;
	 	 	 else if (in >= 395 && in <= 398) out = 2146;
	 	 	 else if (in >= 399 && in <= 402) out = 2147;
	 	 	 else if (in >= 403 && in <= 406) out = 2148;
	 	 	 else if (in >= 407 && in <= 410) out = 2149;
	 	 	 else if (in >= 411 && in <= 414) out = 2150;
	 	 	 else if (in >= 415 && in <= 418) out = 2151;
	 	 	 else if (in >= 419 && in <= 422) out = 2152;
	 	 	 else if (in >= 423 && in <= 426) out = 2153;
	 	 	 else if (in >= 427 && in <= 430) out = 2154;
	 	 	 else if (in >= 431 && in <= 434) out = 2155;
	 	 	 else if (in >= 435 && in <= 438) out = 2156;
	 	 	 else if (in >= 439 && in <= 442) out = 2157;
	 	 	 else if (in >= 443 && in <= 446) out = 2158;
	 	 	 else if (in >= 447 && in <= 450) out = 2159;
	 	 	 else if (in >= 451 && in <= 454) out = 2160;
	 	 	 else if (in >= 455 && in <= 458) out = 2161;
	 	 	 else if (in >= 459 && in <= 462) out = 2162;
	 	 	 else if (in >= 463 && in <= 466) out = 2163;
	 	 	 else if (in >= 467 && in <= 470) out = 2164;
	 	 	 else if (in >= 471 && in <= 474) out = 2165;
	 	 	 else if (in >= 475 && in <= 478) out = 2166;
	 	 	 else if (in >= 479 && in <= 482) out = 2167;
	 	 	 else if (in >= 483 && in <= 486) out = 2168;
	 	 	 else if (in >= 487 && in <= 490) out = 2169;
	 	 	 else if (in >= 491 && in <= 494) out = 2170;
	 	 	 else if (in >= 495 && in <= 498) out = 2171;
	 	 	 else if (in >= 499 && in <= 502) out = 2172;
	 	 	 else if (in >= 503 && in <= 506) out = 2173;
	 	 	 else if (in >= 507 && in <= 510) out = 2174;
	 	 	 else if (in >= 511 && in <= 514) out = 2175;
	 	 	 else if (in >= 515 && in <= 518) out = 2176;
	 	 	 else if (in >= 519 && in <= 522) out = 2177;
	 	 	 else if (in >= 523 && in <= 526) out = 2178;
	 	 	 else if (in >= 527 && in <= 530) out = 2179;
	 	 	 else if (in >= 531 && in <= 534) out = 2180;
	 	 	 else if (in >= 535 && in <= 538) out = 2181;
	 	 	 else if (in >= 539 && in <= 542) out = 2182;
	 	 	 else if (in >= 543 && in <= 546) out = 2183;
	 	 	 else if (in >= 547 && in <= 550) out = 2184;
	 	 	 else if (in >= 551 && in <= 554) out = 2185;
	 	 	 else if (in >= 555 && in <= 559) out = 2186;
	 	 	 else if (in >= 560 && in <= 563) out = 2187;
	 	 	 else if (in >= 564 && in <= 567) out = 2188;
	 	 	 else if (in >= 568 && in <= 571) out = 2189;
	 	 	 else if (in >= 572 && in <= 575) out = 2190;
	 	 	 else if (in >= 576 && in <= 579) out = 2191;
	 	 	 else if (in >= 580 && in <= 583) out = 2192;
	 	 	 else if (in >= 584 && in <= 587) out = 2193;
	 	 	 else if (in >= 588 && in <= 591) out = 2194;
	 	 	 else if (in >= 592 && in <= 595) out = 2195;
	 	 	 else if (in >= 596 && in <= 599) out = 2196;
	 	 	 else if (in >= 600 && in <= 603) out = 2197;
	 	 	 else if (in >= 604 && in <= 607) out = 2198;
	 	 	 else if (in >= 608 && in <= 611) out = 2199;
	 	 	 else if (in >= 612 && in <= 615) out = 2200;
	 	 	 else if (in >= 616 && in <= 619) out = 2201;
	 	 	 else if (in >= 620 && in <= 623) out = 2202;
	 	 	 else if (in >= 624 && in <= 627) out = 2203;
	 	 	 else if (in >= 628 && in <= 631) out = 2204;
	 	 	 else if (in >= 632 && in <= 635) out = 2205;
	 	 	 else if (in >= 636 && in <= 639) out = 2206;
	 	 	 else if (in >= 640 && in <= 643) out = 2207;
	 	 	 else if (in >= 644 && in <= 647) out = 2208;
	 	 	 else if (in >= 648 && in <= 651) out = 2209;
	 	 	 else if (in >= 652 && in <= 655) out = 2210;
	 	 	 else if (in >= 656 && in <= 659) out = 2211;
	 	 	 else if (in >= 660 && in <= 663) out = 2212;
	 	 	 else if (in >= 664 && in <= 667) out = 2213;
	 	 	 else if (in >= 668 && in <= 671) out = 2214;
	 	 	 else if (in >= 672 && in <= 675) out = 2215;
	 	 	 else if (in >= 676 && in <= 679) out = 2216;
	 	 	 else if (in >= 680 && in <= 683) out = 2217;
	 	 	 else if (in >= 684 && in <= 687) out = 2218;
	 	 	 else if (in >= 688 && in <= 691) out = 2219;
	 	 	 else if (in >= 692 && in <= 695) out = 2220;
	 	 	 else if (in >= 696 && in <= 699) out = 2221;
	 	 	 else if (in >= 700 && in <= 703) out = 2222;
	 	 	 else if (in >= 704 && in <= 707) out = 2223;
	 	 	 else if (in >= 708 && in <= 711) out = 2224;
	 	 	 else if (in >= 712 && in <= 715) out = 2225;
	 	 	 else if (in >= 716 && in <= 720) out = 2226;
	 	 	 else if (in >= 721 && in <= 724) out = 2227;
	 	 	 else if (in >= 725 && in <= 728) out = 2228;
	 	 	 else if (in >= 729 && in <= 732) out = 2229;
	 	 	 else if (in >= 733 && in <= 736) out = 2230;
	 	 	 else if (in >= 737 && in <= 740) out = 2231;
	 	 	 else if (in >= 741 && in <= 744) out = 2232;
	 	 	 else if (in >= 745 && in <= 748) out = 2233;
	 	 	 else if (in >= 749 && in <= 752) out = 2234;
	 	 	 else if (in >= 753 && in <= 756) out = 2235;
	 	 	 else if (in >= 757 && in <= 760) out = 2236;
	 	 	 else if (in >= 761 && in <= 764) out = 2237;
	 	 	 else if (in >= 765 && in <= 768) out = 2238;
	 	 	 else if (in >= 769 && in <= 772) out = 2239;
	 	 	 else if (in >= 773 && in <= 776) out = 2240;
	 	 	 else if (in >= 777 && in <= 780) out = 2241;
	 	 	 else if (in >= 781 && in <= 784) out = 2242;
	 	 	 else if (in >= 785 && in <= 788) out = 2243;
	 	 	 else if (in >= 789 && in <= 792) out = 2244;
	 	 	 else if (in >= 793 && in <= 796) out = 2245;
	 	 	 else if (in >= 797 && in <= 800) out = 2246;
	 	 	 else if (in >= 801 && in <= 804) out = 2247;
	 	 	 else if (in >= 805 && in <= 808) out = 2248;
	 	 	 else if (in >= 809 && in <= 812) out = 2249;
	 	 	 else if (in >= 813 && in <= 816) out = 2250;
	 	 	 else if (in >= 817 && in <= 820) out = 2251;
	 	 	 else if (in >= 821 && in <= 824) out = 2252;
	 	 	 else if (in >= 825 && in <= 829) out = 2253;
	 	 	 else if (in >= 830 && in <= 833) out = 2254;
	 	 	 else if (in >= 834 && in <= 837) out = 2255;
	 	 	 else if (in >= 838 && in <= 841) out = 2256;
	 	 	 else if (in >= 842 && in <= 845) out = 2257;
	 	 	 else if (in >= 846 && in <= 849) out = 2258;
	 	 	 else if (in >= 850 && in <= 853) out = 2259;
	 	 	 else if (in >= 854 && in <= 857) out = 2260;
	 	 	 else if (in >= 858 && in <= 861) out = 2261;
	 	 	 else if (in >= 862 && in <= 865) out = 2262;
	 	 	 else if (in >= 866 && in <= 869) out = 2263;
	 	 	 else if (in >= 870 && in <= 873) out = 2264;
	 	 	 else if (in >= 874 && in <= 877) out = 2265;
	 	 	 else if (in >= 878 && in <= 881) out = 2266;
	 	 	 else if (in >= 882 && in <= 885) out = 2267;
	 	 	 else if (in >= 886 && in <= 889) out = 2268;
	 	 	 else if (in >= 890 && in <= 893) out = 2269;
	 	 	 else if (in >= 894 && in <= 897) out = 2270;
	 	 	 else if (in >= 898 && in <= 901) out = 2271;
	 	 	 else if (in >= 902 && in <= 905) out = 2272;
	 	 	 else if (in >= 906 && in <= 909) out = 2273;
	 	 	 else if (in >= 910 && in <= 913) out = 2274;
	 	 	 else if (in >= 914 && in <= 918) out = 2275;
	 	 	 else if (in >= 919 && in <= 922) out = 2276;
	 	 	 else if (in >= 923 && in <= 926) out = 2277;
	 	 	 else if (in >= 927 && in <= 930) out = 2278;
	 	 	 else if (in >= 931 && in <= 934) out = 2279;
	 	 	 else if (in >= 935 && in <= 938) out = 2280;
	 	 	 else if (in >= 939 && in <= 942) out = 2281;
	 	 	 else if (in >= 943 && in <= 946) out = 2282;
	 	 	 else if (in >= 947 && in <= 950) out = 2283;
	 	 	 else if (in >= 951 && in <= 954) out = 2284;
	 	 	 else if (in >= 955 && in <= 958) out = 2285;
	 	 	 else if (in >= 959 && in <= 962) out = 2286;
	 	 	 else if (in >= 963 && in <= 966) out = 2287;
	 	 	 else if (in >= 967 && in <= 970) out = 2288;
	 	 	 else if (in >= 971 && in <= 974) out = 2289;
	 	 	 else if (in >= 975 && in <= 978) out = 2290;
	 	 	 else if (in >= 979 && in <= 982) out = 2291;
	 	 	 else if (in >= 983 && in <= 986) out = 2292;
	 	 	 else if (in >= 987 && in <= 991) out = 2293;
	 	 	 else if (in >= 992 && in <= 995) out = 2294;
	 	 	 else if (in >= 996 && in <= 999) out = 2295;
	 	 	 else if (in >= 1000 && in <= 1003) out = 2296;
	 	 	 else if (in >= 1004 && in <= 1007) out = 2297;
	 	 	 else if (in >= 1008 && in <= 1011) out = 2298;
	 	 	 else if (in >= 1012 && in <= 1015) out = 2299;
	 	 	 else if (in >= 1016 && in <= 1019) out = 2300;
	 	 	 else if (in >= 1020 && in <= 1023) out = 2301;
	 	 	 else if (in >= 1024 && in <= 1027) out = 2302;
	 	 	 else if (in >= 1028 && in <= 1031) out = 2303;
	 	 	 else if (in >= 1032 && in <= 1035) out = 2304;
	 	 	 else if (in >= 1036 && in <= 1039) out = 2305;
	 	 	 else if (in >= 1040 && in <= 1043) out = 2306;
	 	 	 else if (in >= 1044 && in <= 1047) out = 2307;
	 	 	 else if (in >= 1048 && in <= 1052) out = 2308;
	 	 	 else if (in >= 1053 && in <= 1056) out = 2309;
	 	 	 else if (in >= 1057 && in <= 1060) out = 2310;
	 	 	 else if (in >= 1061 && in <= 1064) out = 2311;
	 	 	 else if (in >= 1065 && in <= 1068) out = 2312;
	 	 	 else if (in >= 1069 && in <= 1072) out = 2313;
	 	 	 else if (in >= 1073 && in <= 1076) out = 2314;
	 	 	 else if (in >= 1077 && in <= 1080) out = 2315;
	 	 	 else if (in >= 1081 && in <= 1084) out = 2316;
	 	 	 else if (in >= 1085 && in <= 1088) out = 2317;
	 	 	 else if (in >= 1089 && in <= 1092) out = 2318;
	 	 	 else if (in >= 1093 && in <= 1096) out = 2319;
	 	 	 else if (in >= 1097 && in <= 1100) out = 2320;
	 	 	 else if (in >= 1101 && in <= 1104) out = 2321;
	 	 	 else if (in >= 1105 && in <= 1108) out = 2322;
	 	 	 else if (in >= 1109 && in <= 1113) out = 2323;
	 	 	 else if (in >= 1114 && in <= 1117) out = 2324;
	 	 	 else if (in >= 1118 && in <= 1121) out = 2325;
	 	 	 else if (in >= 1122 && in <= 1125) out = 2326;
	 	 	 else if (in >= 1126 && in <= 1129) out = 2327;
	 	 	 else if (in >= 1130 && in <= 1133) out = 2328;
	 	 	 else if (in >= 1134 && in <= 1137) out = 2329;
	 	 	 else if (in >= 1138 && in <= 1141) out = 2330;
	 	 	 else if (in >= 1142 && in <= 1145) out = 2331;
	 	 	 else if (in >= 1146 && in <= 1149) out = 2332;
	 	 	 else if (in >= 1150 && in <= 1153) out = 2333;
	 	 	 else if (in >= 1154 && in <= 1157) out = 2334;
	 	 	 else if (in >= 1158 && in <= 1162) out = 2335;
	 	 	 else if (in >= 1163 && in <= 1166) out = 2336;
	 	 	 else if (in >= 1167 && in <= 1170) out = 2337;
	 	 	 else if (in >= 1171 && in <= 1174) out = 2338;
	 	 	 else if (in >= 1175 && in <= 1178) out = 2339;
	 	 	 else if (in >= 1179 && in <= 1182) out = 2340;
	 	 	 else if (in >= 1183 && in <= 1186) out = 2341;
	 	 	 else if (in >= 1187 && in <= 1190) out = 2342;
	 	 	 else if (in >= 1191 && in <= 1194) out = 2343;
	 	 	 else if (in >= 1195 && in <= 1198) out = 2344;
	 	 	 else if (in >= 1199 && in <= 1202) out = 2345;
	 	 	 else if (in >= 1203 && in <= 1206) out = 2346;
	 	 	 else if (in >= 1207 && in <= 1211) out = 2347;
	 	 	 else if (in >= 1212 && in <= 1215) out = 2348;
	 	 	 else if (in >= 1216 && in <= 1219) out = 2349;
	 	 	 else if (in >= 1220 && in <= 1223) out = 2350;
	 	 	 else if (in >= 1224 && in <= 1227) out = 2351;
	 	 	 else if (in >= 1228 && in <= 1231) out = 2352;
	 	 	 else if (in >= 1232 && in <= 1235) out = 2353;
	 	 	 else if (in >= 1236 && in <= 1239) out = 2354;
	 	 	 else if (in >= 1240 && in <= 1243) out = 2355;
	 	 	 else if (in >= 1244 && in <= 1247) out = 2356;
	 	 	 else if (in >= 1248 && in <= 1251) out = 2357;
	 	 	 else if (in >= 1252 && in <= 1256) out = 2358;
	 	 	 else if (in >= 1257 && in <= 1260) out = 2359;
	 	 	 else if (in >= 1261 && in <= 1264) out = 2360;
	 	 	 else if (in >= 1265 && in <= 1268) out = 2361;
	 	 	 else if (in >= 1269 && in <= 1272) out = 2362;
	 	 	 else if (in >= 1273 && in <= 1276) out = 2363;
	 	 	 else if (in >= 1277 && in <= 1280) out = 2364;
	 	 	 else if (in >= 1281 && in <= 1284) out = 2365;
	 	 	 else if (in >= 1285 && in <= 1288) out = 2366;
	 	 	 else if (in >= 1289 && in <= 1292) out = 2367;
	 	 	 else if (in >= 1293 && in <= 1297) out = 2368;
	 	 	 else if (in >= 1298 && in <= 1301) out = 2369;
	 	 	 else if (in >= 1302 && in <= 1305) out = 2370;
	 	 	 else if (in >= 1306 && in <= 1309) out = 2371;
	 	 	 else if (in >= 1310 && in <= 1313) out = 2372;
	 	 	 else if (in >= 1314 && in <= 1317) out = 2373;
	 	 	 else if (in >= 1318 && in <= 1321) out = 2374;
	 	 	 else if (in >= 1322 && in <= 1325) out = 2375;
	 	 	 else if (in >= 1326 && in <= 1329) out = 2376;
	 	 	 else if (in >= 1330 && in <= 1333) out = 2377;
	 	 	 else if (in >= 1334 && in <= 1338) out = 2378;
	 	 	 else if (in >= 1339 && in <= 1342) out = 2379;
	 	 	 else if (in >= 1343 && in <= 1346) out = 2380;
	 	 	 else if (in >= 1347 && in <= 1350) out = 2381;
	 	 	 else if (in >= 1351 && in <= 1354) out = 2382;
	 	 	 else if (in >= 1355 && in <= 1358) out = 2383;
	 	 	 else if (in >= 1359 && in <= 1362) out = 2384;
	 	 	 else if (in >= 1363 && in <= 1366) out = 2385;
	 	 	 else if (in >= 1367 && in <= 1370) out = 2386;
	 	 	 else if (in >= 1371 && in <= 1375) out = 2387;
	 	 	 else if (in >= 1376 && in <= 1379) out = 2388;
	 	 	 else if (in >= 1380 && in <= 1383) out = 2389;
	 	 	 else if (in >= 1384 && in <= 1387) out = 2390;
	 	 	 else if (in >= 1388 && in <= 1391) out = 2391;
	 	 	 else if (in >= 1392 && in <= 1395) out = 2392;
	 	 	 else if (in >= 1396 && in <= 1399) out = 2393;
	 	 	 else if (in >= 1400 && in <= 1403) out = 2394;
	 	 	 else if (in >= 1404 && in <= 1408) out = 2395;
	 	 	 else if (in >= 1409 && in <= 1412) out = 2396;
	 	 	 else if (in >= 1413 && in <= 1416) out = 2397;
	 	 	 else if (in >= 1417 && in <= 1420) out = 2398;
	 	 	 else if (in >= 1421 && in <= 1424) out = 2399;
	 	 	 else if (in >= 1425 && in <= 1428) out = 2400;
	 	 	 else if (in >= 1429 && in <= 1432) out = 2401;
	 	 	 else if (in >= 1433 && in <= 1436) out = 2402;
	 	 	 else if (in >= 1437 && in <= 1441) out = 2403;
	 	 	 else if (in >= 1442 && in <= 1445) out = 2404;
	 	 	 else if (in >= 1446 && in <= 1449) out = 2405;
	 	 	 else if (in >= 1450 && in <= 1453) out = 2406;
	 	 	 else if (in >= 1454 && in <= 1457) out = 2407;
	 	 	 else if (in >= 1458 && in <= 1461) out = 2408;
	 	 	 else if (in >= 1462 && in <= 1465) out = 2409;
	 	 	 else if (in >= 1466 && in <= 1469) out = 2410;
	 	 	 else if (in >= 1470 && in <= 1474) out = 2411;
	 	 	 else if (in >= 1475 && in <= 1478) out = 2412;
	 	 	 else if (in >= 1479 && in <= 1482) out = 2413;
	 	 	 else if (in >= 1483 && in <= 1486) out = 2414;
	 	 	 else if (in >= 1487 && in <= 1490) out = 2415;
	 	 	 else if (in >= 1491 && in <= 1494) out = 2416;
	 	 	 else if (in >= 1495 && in <= 1498) out = 2417;
	 	 	 else if (in >= 1499 && in <= 1503) out = 2418;
	 	 	 else if (in >= 1504 && in <= 1507) out = 2419;
	 	 	 else if (in >= 1508 && in <= 1511) out = 2420;
	 	 	 else if (in >= 1512 && in <= 1515) out = 2421;
	 	 	 else if (in >= 1516 && in <= 1519) out = 2422;
	 	 	 else if (in >= 1520 && in <= 1523) out = 2423;
	 	 	 else if (in >= 1524 && in <= 1527) out = 2424;
	 	 	 else if (in >= 1528 && in <= 1531) out = 2425;
	 	 	 else if (in >= 1532 && in <= 1536) out = 2426;
	 	 	 else if (in >= 1537 && in <= 1540) out = 2427;
	 	 	 else if (in >= 1541 && in <= 1544) out = 2428;
	 	 	 else if (in >= 1545 && in <= 1548) out = 2429;
	 	 	 else if (in >= 1549 && in <= 1552) out = 2430;
	 	 	 else if (in >= 1553 && in <= 1556) out = 2431;
	 	 	 else if (in >= 1557 && in <= 1560) out = 2432;
	 	 	 else if (in >= 1561 && in <= 1565) out = 2433;
	 	 	 else if (in >= 1566 && in <= 1569) out = 2434;
	 	 	 else if (in >= 1570 && in <= 1573) out = 2435;
	 	 	 else if (in >= 1574 && in <= 1577) out = 2436;
	 	 	 else if (in >= 1578 && in <= 1581) out = 2437;
	 	 	 else if (in >= 1582 && in <= 1585) out = 2438;
	 	 	 else if (in >= 1586 && in <= 1590) out = 2439;
	 	 	 else if (in >= 1591 && in <= 1594) out = 2440;
	 	 	 else if (in >= 1595 && in <= 1598) out = 2441;
	 	 	 else if (in >= 1599 && in <= 1602) out = 2442;
	 	 	 else if (in >= 1603 && in <= 1606) out = 2443;
	 	 	 else if (in >= 1607 && in <= 1610) out = 2444;
	 	 	 else if (in >= 1611 && in <= 1614) out = 2445;
	 	 	 else if (in >= 1615 && in <= 1619) out = 2446;
	 	 	 else if (in >= 1620 && in <= 1623) out = 2447;
	 	 	 else if (in >= 1624 && in <= 1627) out = 2448;
	 	 	 else if (in >= 1628 && in <= 1631) out = 2449;
	 	 	 else if (in >= 1632 && in <= 1635) out = 2450;
	 	 	 else if (in >= 1636 && in <= 1639) out = 2451;
	 	 	 else if (in >= 1640 && in <= 1644) out = 2452;
	 	 	 else if (in >= 1645 && in <= 1648) out = 2453;
	 	 	 else if (in >= 1649 && in <= 1652) out = 2454;
	 	 	 else if (in >= 1653 && in <= 1656) out = 2455;
	 	 	 else if (in >= 1657 && in <= 1660) out = 2456;
	 	 	 else if (in >= 1661 && in <= 1664) out = 2457;
	 	 	 else if (in >= 1665 && in <= 1669) out = 2458;
	 	 	 else if (in >= 1670 && in <= 1673) out = 2459;
	 	 	 else if (in >= 1674 && in <= 1677) out = 2460;
	 	 	 else if (in >= 1678 && in <= 1681) out = 2461;
	 	 	 else if (in >= 1682 && in <= 1685) out = 2462;
	 	 	 else if (in >= 1686 && in <= 1689) out = 2463;
	 	 	 else if (in >= 1690 && in <= 1694) out = 2464;
	 	 	 else if (in >= 1695 && in <= 1698) out = 2465;
	 	 	 else if (in >= 1699 && in <= 1702) out = 2466;
	 	 	 else if (in >= 1703 && in <= 1706) out = 2467;
	 	 	 else if (in >= 1707 && in <= 1710) out = 2468;
	 	 	 else if (in >= 1711 && in <= 1715) out = 2469;
	 	 	 else if (in >= 1716 && in <= 1719) out = 2470;
	 	 	 else if (in >= 1720 && in <= 1723) out = 2471;
	 	 	 else if (in >= 1724 && in <= 1727) out = 2472;
	 	 	 else if (in >= 1728 && in <= 1731) out = 2473;
	 	 	 else if (in >= 1732 && in <= 1735) out = 2474;
	 	 	 else if (in >= 1736 && in <= 1740) out = 2475;
	 	 	 else if (in >= 1741 && in <= 1744) out = 2476;
	 	 	 else if (in >= 1745 && in <= 1748) out = 2477;
	 	 	 else if (in >= 1749 && in <= 1752) out = 2478;
	 	 	 else if (in >= 1753 && in <= 1756) out = 2479;
	 	 	 else if (in >= 1757 && in <= 1761) out = 2480;
	 	 	 else if (in >= 1762 && in <= 1765) out = 2481;
	 	 	 else if (in >= 1766 && in <= 1769) out = 2482;
	 	 	 else if (in >= 1770 && in <= 1773) out = 2483;
	 	 	 else if (in >= 1774 && in <= 1777) out = 2484;
	 	 	 else if (in >= 1778 && in <= 1782) out = 2485;
	 	 	 else if (in >= 1783 && in <= 1786) out = 2486;
	 	 	 else if (in >= 1787 && in <= 1790) out = 2487;
	 	 	 else if (in >= 1791 && in <= 1794) out = 2488;
	 	 	 else if (in >= 1795 && in <= 1798) out = 2489;
	 	 	 else if (in >= 1799 && in <= 1802) out = 2490;
	 	 	 else if (in >= 1803 && in <= 1807) out = 2491;
	 	 	 else if (in >= 1808 && in <= 1811) out = 2492;
	 	 	 else if (in >= 1812 && in <= 1815) out = 2493;
	 	 	 else if (in >= 1816 && in <= 1819) out = 2494;
	 	 	 else if (in >= 1820 && in <= 1823) out = 2495;
	 	 	 else if (in >= 1824 && in <= 1828) out = 2496;
	 	 	 else if (in >= 1829 && in <= 1832) out = 2497;
	 	 	 else if (in >= 1833 && in <= 1836) out = 2498;
	 	 	 else if (in >= 1837 && in <= 1840) out = 2499;
	 	 	 else if (in >= 1841 && in <= 1845) out = 2500;
	 	 	 else if (in >= 1846 && in <= 1849) out = 2501;
	 	 	 else if (in >= 1850 && in <= 1853) out = 2502;
	 	 	 else if (in >= 1854 && in <= 1857) out = 2503;
	 	 	 else if (in >= 1858 && in <= 1861) out = 2504;
	 	 	 else if (in >= 1862 && in <= 1866) out = 2505;
	 	 	 else if (in >= 1867 && in <= 1870) out = 2506;
	 	 	 else if (in >= 1871 && in <= 1874) out = 2507;
	 	 	 else if (in >= 1875 && in <= 1878) out = 2508;
	 	 	 else if (in >= 1879 && in <= 1882) out = 2509;
	 	 	 else if (in >= 1883 && in <= 1887) out = 2510;
	 	 	 else if (in >= 1888 && in <= 1891) out = 2511;
	 	 	 else if (in >= 1892 && in <= 1895) out = 2512;
	 	 	 else if (in >= 1896 && in <= 1899) out = 2513;
	 	 	 else if (in >= 1900 && in <= 1904) out = 2514;
	 	 	 else if (in >= 1905 && in <= 1908) out = 2515;
	 	 	 else if (in >= 1909 && in <= 1912) out = 2516;
	 	 	 else if (in >= 1913 && in <= 1916) out = 2517;
	 	 	 else if (in >= 1917 && in <= 1920) out = 2518;
	 	 	 else if (in >= 1921 && in <= 1925) out = 2519;
	 	 	 else if (in >= 1926 && in <= 1929) out = 2520;
	 	 	 else if (in >= 1930 && in <= 1933) out = 2521;
	 	 	 else if (in >= 1934 && in <= 1937) out = 2522;
	 	 	 else if (in >= 1938 && in <= 1942) out = 2523;
	 	 	 else if (in >= 1943 && in <= 1946) out = 2524;
	 	 	 else if (in >= 1947 && in <= 1950) out = 2525;
	 	 	 else if (in >= 1951 && in <= 1954) out = 2526;
	 	 	 else if (in >= 1955 && in <= 1958) out = 2527;
	 	 	 else if (in >= 1959 && in <= 1963) out = 2528;
	 	 	 else if (in >= 1964 && in <= 1967) out = 2529;
	 	 	 else if (in >= 1968 && in <= 1971) out = 2530;
	 	 	 else if (in >= 1972 && in <= 1975) out = 2531;
	 	 	 else if (in >= 1976 && in <= 1980) out = 2532;
	 	 	 else if (in >= 1981 && in <= 1984) out = 2533;
	 	 	 else if (in >= 1985 && in <= 1988) out = 2534;
	 	 	 else if (in >= 1989 && in <= 1992) out = 2535;
	 	 	 else if (in >= 1993 && in <= 1997) out = 2536;
	 	 	 else if (in >= 1998 && in <= 2001) out = 2537;
	 	 	 else if (in >= 2002 && in <= 2005) out = 2538;
	 	 	 else if (in >= 2006 && in <= 2009) out = 2539;
	 	 	 else if (in >= 2010 && in <= 2014) out = 2540;
	 	 	 else if (in >= 2015 && in <= 2018) out = 2541;
	 	 	 else if (in >= 2019 && in <= 2022) out = 2542;
	 	 	 else if (in >= 2023 && in <= 2026) out = 2543;
	 	 	 else if (in >= 2027 && in <= 2031) out = 2544;
	 	 	 else if (in >= 2032 && in <= 2035) out = 2545;
	 	 	 else if (in >= 2036 && in <= 2039) out = 2546;
	 	 	 else if (in >= 2040 && in <= 2043) out = 2547;
	 	 	 else if (in >= 2044 && in <= 2048) out = 2548;
	 	 	 else if (in >= 2049 && in <= 2052) out = 2549;
	 	 	 else if (in >= 2053 && in <= 2056) out = 2550;
	 	 	 else if (in >= 2057 && in <= 2060) out = 2551;
	 	 	 else if (in >= 2061 && in <= 2065) out = 2552;
	 	 	 else if (in >= 2066 && in <= 2069) out = 2553;
	 	 	 else if (in >= 2070 && in <= 2073) out = 2554;
	 	 	 else if (in >= 2074 && in <= 2077) out = 2555;
	 	 	 else if (in >= 2078 && in <= 2082) out = 2556;
	 	 	 else if (in >= 2083 && in <= 2086) out = 2557;
	 	 	 else if (in >= 2087 && in <= 2090) out = 2558;
	 	 	 else if (in >= 2091 && in <= 2095) out = 2559;
	 	 	 else if (in >= 2096 && in <= 2099) out = 2560;
	 	 	 else if (in >= 2100 && in <= 2103) out = 2561;
	 	 	 else if (in >= 2104 && in <= 2107) out = 2562;
	 	 	 else if (in >= 2108 && in <= 2112) out = 2563;
	 	 	 else if (in >= 2113 && in <= 2116) out = 2564;
	 	 	 else if (in >= 2117 && in <= 2120) out = 2565;
	 	 	 else if (in >= 2121 && in <= 2124) out = 2566;
	 	 	 else if (in >= 2125 && in <= 2129) out = 2567;
	 	 	 else if (in >= 2130 && in <= 2133) out = 2568;
	 	 	 else if (in >= 2134 && in <= 2137) out = 2569;
	 	 	 else if (in >= 2138 && in <= 2142) out = 2570;
	 	 	 else if (in >= 2143 && in <= 2146) out = 2571;
	 	 	 else if (in >= 2147 && in <= 2150) out = 2572;
	 	 	 else if (in >= 2151 && in <= 2154) out = 2573;
	 	 	 else if (in >= 2155 && in <= 2159) out = 2574;
	 	 	 else if (in >= 2160 && in <= 2163) out = 2575;
	 	 	 else if (in >= 2164 && in <= 2167) out = 2576;
	 	 	 else if (in >= 2168 && in <= 2172) out = 2577;
	 	 	 else if (in >= 2173 && in <= 2176) out = 2578;
	 	 	 else if (in >= 2177 && in <= 2180) out = 2579;
	 	 	 else if (in >= 2181 && in <= 2184) out = 2580;
	 	 	 else if (in >= 2185 && in <= 2189) out = 2581;
	 	 	 else if (in >= 2190 && in <= 2193) out = 2582;
	 	 	 else if (in >= 2194 && in <= 2197) out = 2583;
	 	 	 else if (in >= 2198 && in <= 2202) out = 2584;
	 	 	 else if (in >= 2203 && in <= 2206) out = 2585;
	 	 	 else if (in >= 2207 && in <= 2210) out = 2586;
	 	 	 else if (in >= 2211 && in <= 2214) out = 2587;
	 	 	 else if (in >= 2215 && in <= 2219) out = 2588;
	 	 	 else if (in >= 2220 && in <= 2223) out = 2589;
	 	 	 else if (in >= 2224 && in <= 2227) out = 2590;
	 	 	 else if (in >= 2228 && in <= 2232) out = 2591;
	 	 	 else if (in >= 2233 && in <= 2236) out = 2592;
	 	 	 else if (in >= 2237 && in <= 2240) out = 2593;
	 	 	 else if (in >= 2241 && in <= 2245) out = 2594;
	 	 	 else if (in >= 2246 && in <= 2249) out = 2595;
	 	 	 else if (in >= 2250 && in <= 2253) out = 2596;
	 	 	 else if (in >= 2254 && in <= 2258) out = 2597;
	 	 	 else if (in >= 2259 && in <= 2262) out = 2598;
	 	 	 else if (in >= 2263 && in <= 2266) out = 2599;
	 	 	 else if (in >= 2267 && in <= 2270) out = 2600;
	 	 	 else if (in >= 2271 && in <= 2275) out = 2601;
	 	 	 else if (in >= 2276 && in <= 2279) out = 2602;
	 	 	 else if (in >= 2280 && in <= 2283) out = 2603;
	 	 	 else if (in >= 2284 && in <= 2288) out = 2604;
	 	 	 else if (in >= 2289 && in <= 2292) out = 2605;
	 	 	 else if (in >= 2293 && in <= 2296) out = 2606;
	 	 	 else if (in >= 2297 && in <= 2301) out = 2607;
	 	 	 else if (in >= 2302 && in <= 2305) out = 2608;
	 	 	 else if (in >= 2306 && in <= 2309) out = 2609;
	 	 	 else if (in >= 2310 && in <= 2314) out = 2610;
	 	 	 else if (in >= 2315 && in <= 2318) out = 2611;
	 	 	 else if (in >= 2319 && in <= 2322) out = 2612;
	 	 	 else if (in >= 2323 && in <= 2327) out = 2613;
	 	 	 else if (in >= 2328 && in <= 2331) out = 2614;
	 	 	 else if (in >= 2332 && in <= 2335) out = 2615;
	 	 	 else if (in >= 2336 && in <= 2340) out = 2616;
	 	 	 else if (in >= 2341 && in <= 2344) out = 2617;
	 	 	 else if (in >= 2345 && in <= 2348) out = 2618;
	 	 	 else if (in >= 2349 && in <= 2353) out = 2619;
	 	 	 else if (in >= 2354 && in <= 2357) out = 2620;
	 	 	 else if (in >= 2358 && in <= 2361) out = 2621;
	 	 	 else if (in >= 2362 && in <= 2366) out = 2622;
	 	 	 else if (in >= 2367 && in <= 2370) out = 2623;
	 	 	 else if (in >= 2371 && in <= 2374) out = 2624;
	 	 	 else if (in >= 2375 && in <= 2379) out = 2625;
	 	 	 else if (in >= 2380 && in <= 2383) out = 2626;
	 	 	 else if (in >= 2384 && in <= 2387) out = 2627;
	 	 	 else if (in >= 2388 && in <= 2392) out = 2628;
	 	 	 else if (in >= 2393 && in <= 2396) out = 2629;
	 	 	 else if (in >= 2397 && in <= 2401) out = 2630;
	 	 	 else if (in >= 2402 && in <= 2405) out = 2631;
	 	 	 else if (in >= 2406 && in <= 2409) out = 2632;
	 	 	 else if (in >= 2410 && in <= 2414) out = 2633;
	 	 	 else if (in >= 2415 && in <= 2418) out = 2634;
	 	 	 else if (in >= 2419 && in <= 2422) out = 2635;
	 	 	 else if (in >= 2423 && in <= 2427) out = 2636;
	 	 	 else if (in >= 2428 && in <= 2431) out = 2637;
	 	 	 else if (in >= 2432 && in <= 2435) out = 2638;
	 	 	 else if (in >= 2436 && in <= 2440) out = 2639;
	 	 	 else if (in >= 2441 && in <= 2444) out = 2640;
	 	 	 else if (in >= 2445 && in <= 2449) out = 2641;
	 	 	 else if (in >= 2450 && in <= 2453) out = 2642;
	 	 	 else if (in >= 2454 && in <= 2457) out = 2643;
	 	 	 else if (in >= 2458 && in <= 2462) out = 2644;
	 	 	 else if (in >= 2463 && in <= 2466) out = 2645;
	 	 	 else if (in >= 2467 && in <= 2470) out = 2646;
	 	 	 else if (in >= 2471 && in <= 2475) out = 2647;
	 	 	 else if (in >= 2476 && in <= 2479) out = 2648;
	 	 	 else if (in >= 2480 && in <= 2484) out = 2649;
	 	 	 else if (in >= 2485 && in <= 2488) out = 2650;
	 	 	 else if (in >= 2489 && in <= 2492) out = 2651;
	 	 	 else if (in >= 2493 && in <= 2497) out = 2652;
	 	 	 else if (in >= 2498 && in <= 2501) out = 2653;
	 	 	 else if (in >= 2502 && in <= 2505) out = 2654;
	 	 	 else if (in >= 2506 && in <= 2510) out = 2655;
	 	 	 else if (in >= 2511 && in <= 2514) out = 2656;
	 	 	 else if (in >= 2515 && in <= 2519) out = 2657;
	 	 	 else if (in >= 2520 && in <= 2523) out = 2658;
	 	 	 else if (in >= 2524 && in <= 2527) out = 2659;
	 	 	 else if (in >= 2528 && in <= 2532) out = 2660;
	 	 	 else if (in >= 2533 && in <= 2536) out = 2661;
	 	 	 else if (in >= 2537 && in <= 2541) out = 2662;
	 	 	 else if (in >= 2542 && in <= 2545) out = 2663;
	 	 	 else if (in >= 2546 && in <= 2549) out = 2664;
	 	 	 else if (in >= 2550 && in <= 2554) out = 2665;
	 	 	 else if (in >= 2555 && in <= 2558) out = 2666;
	 	 	 else if (in >= 2559 && in <= 2563) out = 2667;
	 	 	 else if (in >= 2564 && in <= 2567) out = 2668;
	 	 	 else if (in >= 2568 && in <= 2571) out = 2669;
	 	 	 else if (in >= 2572 && in <= 2576) out = 2670;
	 	 	 else if (in >= 2577 && in <= 2580) out = 2671;
	 	 	 else if (in >= 2581 && in <= 2585) out = 2672;
	 	 	 else if (in >= 2586 && in <= 2589) out = 2673;
	 	 	 else if (in >= 2590 && in <= 2593) out = 2674;
	 	 	 else if (in >= 2594 && in <= 2598) out = 2675;
	 	 	 else if (in >= 2599 && in <= 2602) out = 2676;
	 	 	 else if (in >= 2603 && in <= 2607) out = 2677;
	 	 	 else if (in >= 2608 && in <= 2611) out = 2678;
	 	 	 else if (in >= 2612 && in <= 2616) out = 2679;
	 	 	 else if (in >= 2617 && in <= 2620) out = 2680;
	 	 	 else if (in >= 2621 && in <= 2624) out = 2681;
	 	 	 else if (in >= 2625 && in <= 2629) out = 2682;
	 	 	 else if (in >= 2630 && in <= 2633) out = 2683;
	 	 	 else if (in >= 2634 && in <= 2638) out = 2684;
	 	 	 else if (in >= 2639 && in <= 2642) out = 2685;
	 	 	 else if (in >= 2643 && in <= 2647) out = 2686;
	 	 	 else if (in >= 2648 && in <= 2651) out = 2687;
	 	 	 else if (in >= 2652 && in <= 2655) out = 2688;
	 	 	 else if (in >= 2656 && in <= 2660) out = 2689;
	 	 	 else if (in >= 2661 && in <= 2664) out = 2690;
	 	 	 else if (in >= 2665 && in <= 2669) out = 2691;
	 	 	 else if (in >= 2670 && in <= 2673) out = 2692;
	 	 	 else if (in >= 2674 && in <= 2678) out = 2693;
	 	 	 else if (in >= 2679 && in <= 2682) out = 2694;
	 	 	 else if (in >= 2683 && in <= 2687) out = 2695;
	 	 	 else if (in >= 2688 && in <= 2691) out = 2696;
	 	 	 else if (in >= 2692 && in <= 2695) out = 2697;
	 	 	 else if (in >= 2696 && in <= 2700) out = 2698;
	 	 	 else if (in >= 2701 && in <= 2704) out = 2699;
	 	 	 else if (in >= 2705 && in <= 2709) out = 2700;
	 	 	 else if (in >= 2710 && in <= 2713) out = 2701;
	 	 	 else if (in >= 2714 && in <= 2718) out = 2702;
	 	 	 else if (in >= 2719 && in <= 2722) out = 2703;
	 	 	 else if (in >= 2723 && in <= 2727) out = 2704;
	 	 	 else if (in >= 2728 && in <= 2731) out = 2705;
	 	 	 else if (in >= 2732 && in <= 2736) out = 2706;
	 	 	 else if (in >= 2737 && in <= 2740) out = 2707;
	 	 	 else if (in >= 2741 && in <= 2744) out = 2708;
	 	 	 else if (in >= 2745 && in <= 2749) out = 2709;
	 	 	 else if (in >= 2750 && in <= 2753) out = 2710;
	 	 	 else if (in >= 2754 && in <= 2758) out = 2711;
	 	 	 else if (in >= 2759 && in <= 2762) out = 2712;
	 	 	 else if (in >= 2763 && in <= 2767) out = 2713;
	 	 	 else if (in >= 2768 && in <= 2771) out = 2714;
	 	 	 else if (in >= 2772 && in <= 2776) out = 2715;
	 	 	 else if (in >= 2777 && in <= 2780) out = 2716;
	 	 	 else if (in >= 2781 && in <= 2785) out = 2717;
	 	 	 else if (in >= 2786 && in <= 2789) out = 2718;
	 	 	 else if (in >= 2790 && in <= 2794) out = 2719;
	 	 	 else if (in >= 2795 && in <= 2798) out = 2720;
	 	 	 else if (in >= 2799 && in <= 2803) out = 2721;
	 	 	 else if (in >= 2804 && in <= 2807) out = 2722;
	 	 	 else if (in >= 2808 && in <= 2812) out = 2723;
	 	 	 else if (in >= 2813 && in <= 2816) out = 2724;
	 	 	 else if (in >= 2817 && in <= 2821) out = 2725;
	 	 	 else if (in >= 2822 && in <= 2825) out = 2726;
	 	 	 else if (in >= 2826 && in <= 2830) out = 2727;
	 	 	 else if (in >= 2831 && in <= 2834) out = 2728;
	 	 	 else if (in >= 2835 && in <= 2839) out = 2729;
	 	 	 else if (in >= 2840 && in <= 2843) out = 2730;
	 	 	 else if (in >= 2844 && in <= 2848) out = 2731;
	 	 	 else if (in >= 2849 && in <= 2852) out = 2732;
	 	 	 else if (in >= 2853 && in <= 2857) out = 2733;
	 	 	 else if (in >= 2858 && in <= 2861) out = 2734;
	 	 	 else if (in >= 2862 && in <= 2866) out = 2735;
	 	 	 else if (in >= 2867 && in <= 2870) out = 2736;
	 	 	 else if (in >= 2871 && in <= 2875) out = 2737;
	 	 	 else if (in >= 2876 && in <= 2879) out = 2738;
	 	 	 else if (in >= 2880 && in <= 2884) out = 2739;
	 	 	 else if (in >= 2885 && in <= 2888) out = 2740;
	 	 	 else if (in >= 2889 && in <= 2893) out = 2741;
	 	 	 else if (in >= 2894 && in <= 2897) out = 2742;
	 	 	 else if (in >= 2898 && in <= 2902) out = 2743;
	 	 	 else if (in >= 2903 && in <= 2906) out = 2744;
	 	 	 else if (in >= 2907 && in <= 2911) out = 2745;
	 	 	 else if (in >= 2912 && in <= 2915) out = 2746;
	 	 	 else if (in >= 2916 && in <= 2920) out = 2747;
	 	 	 else if (in >= 2921 && in <= 2924) out = 2748;
	 	 	 else if (in >= 2925 && in <= 2929) out = 2749;
	 	 	 else if (in >= 2930 && in <= 2934) out = 2750;
	 	 	 else if (in >= 2935 && in <= 2938) out = 2751;
	 	 	 else if (in >= 2939 && in <= 2943) out = 2752;
	 	 	 else if (in >= 2944 && in <= 2947) out = 2753;
	 	 	 else if (in >= 2948 && in <= 2952) out = 2754;
	 	 	 else if (in >= 2953 && in <= 2956) out = 2755;
	 	 	 else if (in >= 2957 && in <= 2961) out = 2756;
	 	 	 else if (in >= 2962 && in <= 2965) out = 2757;
	 	 	 else if (in >= 2966 && in <= 2970) out = 2758;
	 	 	 else if (in >= 2971 && in <= 2974) out = 2759;
	 	 	 else if (in >= 2975 && in <= 2979) out = 2760;
	 	 	 else if (in >= 2980 && in <= 2984) out = 2761;
	 	 	 else if (in >= 2985 && in <= 2988) out = 2762;
	 	 	 else if (in >= 2989 && in <= 2993) out = 2763;
	 	 	 else if (in >= 2994 && in <= 2997) out = 2764;
	 	 	 else if (in >= 2998 && in <= 3002) out = 2765;
	 	 	 else if (in >= 3003 && in <= 3006) out = 2766;
	 	 	 else if (in >= 3007 && in <= 3011) out = 2767;
	 	 	 else if (in >= 3012 && in <= 3015) out = 2768;
	 	 	 else if (in >= 3016 && in <= 3020) out = 2769;
	 	 	 else if (in >= 3021 && in <= 3025) out = 2770;
	 	 	 else if (in >= 3026 && in <= 3029) out = 2771;
	 	 	 else if (in >= 3030 && in <= 3034) out = 2772;
	 	 	 else if (in >= 3035 && in <= 3038) out = 2773;
	 	 	 else if (in >= 3039 && in <= 3043) out = 2774;
	 	 	 else if (in >= 3044 && in <= 3047) out = 2775;
	 	 	 else if (in >= 3048 && in <= 3052) out = 2776;
	 	 	 else if (in >= 3053 && in <= 3057) out = 2777;
	 	 	 else if (in >= 3058 && in <= 3061) out = 2778;
	 	 	 else if (in >= 3062 && in <= 3066) out = 2779;
	 	 	 else if (in >= 3067 && in <= 3070) out = 2780;
	 	 	 else if (in >= 3071 && in <= 3075) out = 2781;
	 	 	 else if (in >= 3076 && in <= 3080) out = 2782;
	 	 	 else if (in >= 3081 && in <= 3084) out = 2783;
	 	 	 else if (in >= 3085 && in <= 3089) out = 2784;
	 	 	 else if (in >= 3090 && in <= 3093) out = 2785;
	 	 	 else if (in >= 3094 && in <= 3098) out = 2786;
	 	 	 else if (in >= 3099 && in <= 3103) out = 2787;
	 	 	 else if (in >= 3104 && in <= 3107) out = 2788;
	 	 	 else if (in >= 3108 && in <= 3112) out = 2789;
	 	 	 else if (in >= 3113 && in <= 3116) out = 2790;
	 	 	 else if (in >= 3117 && in <= 3121) out = 2791;
	 	 	 else if (in >= 3122 && in <= 3126) out = 2792;
	 	 	 else if (in >= 3127 && in <= 3130) out = 2793;
	 	 	 else if (in >= 3131 && in <= 3135) out = 2794;
	 	 	 else if (in >= 3136 && in <= 3139) out = 2795;
	 	 	 else if (in >= 3140 && in <= 3144) out = 2796;
	 	 	 else if (in >= 3145 && in <= 3149) out = 2797;
	 	 	 else if (in >= 3150 && in <= 3153) out = 2798;
	 	 	 else if (in >= 3154 && in <= 3158) out = 2799;
	 	 	 else if (in >= 3159 && in <= 3163) out = 2800;
	 	 	 else if (in >= 3164 && in <= 3167) out = 2801;
	 	 	 else if (in >= 3168 && in <= 3172) out = 2802;
	 	 	 else if (in >= 3173 && in <= 3176) out = 2803;
	 	 	 else if (in >= 3177 && in <= 3181) out = 2804;
	 	 	 else if (in >= 3182 && in <= 3186) out = 2805;
	 	 	 else if (in >= 3187 && in <= 3190) out = 2806;
	 	 	 else if (in >= 3191 && in <= 3195) out = 2807;
	 	 	 else if (in >= 3196 && in <= 3200) out = 2808;
	 	 	 else if (in >= 3201 && in <= 3204) out = 2809;
	 	 	 else if (in >= 3205 && in <= 3209) out = 2810;
	 	 	 else if (in >= 3210 && in <= 3214) out = 2811;
	 	 	 else if (in >= 3215 && in <= 3218) out = 2812;
	 	 	 else if (in >= 3219 && in <= 3223) out = 2813;
	 	 	 else if (in >= 3224 && in <= 3228) out = 2814;
	 	 	 else if (in >= 3229 && in <= 3232) out = 2815;
	 	 	 else if (in >= 3233 && in <= 3237) out = 2816;
	 	 	 else if (in >= 3238 && in <= 3242) out = 2817;
	 	 	 else if (in >= 3243 && in <= 3246) out = 2818;
	 	 	 else if (in >= 3247 && in <= 3251) out = 2819;
	 	 	 else if (in >= 3252 && in <= 3256) out = 2820;
	 	 	 else if (in >= 3257 && in <= 3260) out = 2821;
	 	 	 else if (in >= 3261 && in <= 3265) out = 2822;
	 	 	 else if (in >= 3266 && in <= 3270) out = 2823;
	 	 	 else if (in >= 3271 && in <= 3274) out = 2824;
	 	 	 else if (in >= 3275 && in <= 3279) out = 2825;
	 	 	 else if (in >= 3280 && in <= 3284) out = 2826;
	 	 	 else if (in >= 3285 && in <= 3288) out = 2827;
	 	 	 else if (in >= 3289 && in <= 3293) out = 2828;
	 	 	 else if (in >= 3294 && in <= 3298) out = 2829;
	 	 	 else if (in >= 3299 && in <= 3302) out = 2830;
	 	 	 else if (in >= 3303 && in <= 3307) out = 2831;
	 	 	 else if (in >= 3308 && in <= 3312) out = 2832;
	 	 	 else if (in >= 3313 && in <= 3316) out = 2833;
	 	 	 else if (in >= 3317 && in <= 3321) out = 2834;
	 	 	 else if (in >= 3322 && in <= 3326) out = 2835;
	 	 	 else if (in >= 3327 && in <= 3330) out = 2836;
	 	 	 else if (in >= 3331 && in <= 3335) out = 2837;
	 	 	 else if (in >= 3336 && in <= 3340) out = 2838;
	 	 	 else if (in >= 3341 && in <= 3345) out = 2839;
	 	 	 else if (in >= 3346 && in <= 3349) out = 2840;
	 	 	 else if (in >= 3350 && in <= 3354) out = 2841;
	 	 	 else if (in >= 3355 && in <= 3359) out = 2842;
	 	 	 else if (in >= 3360 && in <= 3363) out = 2843;
	 	 	 else if (in >= 3364 && in <= 3368) out = 2844;
	 	 	 else if (in >= 3369 && in <= 3373) out = 2845;
	 	 	 else if (in >= 3374 && in <= 3378) out = 2846;
	 	 	 else if (in >= 3379 && in <= 3382) out = 2847;
	 	 	 else if (in >= 3383 && in <= 3387) out = 2848;
	 	 	 else if (in >= 3388 && in <= 3392) out = 2849;
	 	 	 else if (in >= 3393 && in <= 3396) out = 2850;
	 	 	 else if (in >= 3397 && in <= 3401) out = 2851;
	 	 	 else if (in >= 3402 && in <= 3406) out = 2852;
	 	 	 else if (in >= 3407 && in <= 3411) out = 2853;
	 	 	 else if (in >= 3412 && in <= 3415) out = 2854;
	 	 	 else if (in >= 3416 && in <= 3420) out = 2855;
	 	 	 else if (in >= 3421 && in <= 3425) out = 2856;
	 	 	 else if (in >= 3426 && in <= 3430) out = 2857;
	 	 	 else if (in >= 3431 && in <= 3434) out = 2858;
	 	 	 else if (in >= 3435 && in <= 3439) out = 2859;
	 	 	 else if (in >= 3440 && in <= 3444) out = 2860;
	 	 	 else if (in >= 3445 && in <= 3449) out = 2861;
	 	 	 else if (in >= 3450 && in <= 3453) out = 2862;
	 	 	 else if (in >= 3454 && in <= 3458) out = 2863;
	 	 	 else if (in >= 3459 && in <= 3463) out = 2864;
	 	 	 else if (in >= 3464 && in <= 3468) out = 2865;
	 	 	 else if (in >= 3469 && in <= 3472) out = 2866;
	 	 	 else if (in >= 3473 && in <= 3477) out = 2867;
	 	 	 else if (in >= 3478 && in <= 3482) out = 2868;
	 	 	 else if (in >= 3483 && in <= 3487) out = 2869;
	 	 	 else if (in >= 3488 && in <= 3491) out = 2870;
	 	 	 else if (in >= 3492 && in <= 3496) out = 2871;
	 	 	 else if (in >= 3497 && in <= 3501) out = 2872;
	 	 	 else if (in >= 3502 && in <= 3506) out = 2873;
	 	 	 else if (in >= 3507 && in <= 3511) out = 2874;
	 	 	 else if (in >= 3512 && in <= 3515) out = 2875;
	 	 	 else if (in >= 3516 && in <= 3520) out = 2876;
	 	 	 else if (in >= 3521 && in <= 3525) out = 2877;
	 	 	 else if (in >= 3526 && in <= 3530) out = 2878;
	 	 	 else if (in >= 3531 && in <= 3535) out = 2879;
	 	 	 else if (in >= 3536 && in <= 3539) out = 2880;
	 	 	 else if (in >= 3540 && in <= 3544) out = 2881;
	 	 	 else if (in >= 3545 && in <= 3549) out = 2882;
	 	 	 else if (in >= 3550 && in <= 3554) out = 2883;
	 	 	 else if (in >= 3555 && in <= 3559) out = 2884;
	 	 	 else if (in >= 3560 && in <= 3563) out = 2885;
	 	 	 else if (in >= 3564 && in <= 3568) out = 2886;
	 	 	 else if (in >= 3569 && in <= 3573) out = 2887;
	 	 	 else if (in >= 3574 && in <= 3578) out = 2888;
	 	 	 else if (in >= 3579 && in <= 3583) out = 2889;
	 	 	 else if (in >= 3584 && in <= 3587) out = 2890;
	 	 	 else if (in >= 3588 && in <= 3592) out = 2891;
	 	 	 else if (in >= 3593 && in <= 3597) out = 2892;
	 	 	 else if (in >= 3598 && in <= 3602) out = 2893;
	 	 	 else if (in >= 3603 && in <= 3607) out = 2894;
	 	 	 else if (in >= 3608 && in <= 3612) out = 2895;
	 	 	 else if (in >= 3613 && in <= 3616) out = 2896;
	 	 	 else if (in >= 3617 && in <= 3621) out = 2897;
	 	 	 else if (in >= 3622 && in <= 3626) out = 2898;
	 	 	 else if (in >= 3627 && in <= 3631) out = 2899;
	 	 	 else if (in >= 3632 && in <= 3636) out = 2900;
	 	 	 else if (in >= 3637 && in <= 3641) out = 2901;
	 	 	 else if (in >= 3642 && in <= 3645) out = 2902;
	 	 	 else if (in >= 3646 && in <= 3650) out = 2903;
	 	 	 else if (in >= 3651 && in <= 3655) out = 2904;
	 	 	 else if (in >= 3656 && in <= 3660) out = 2905;
	 	 	 else if (in >= 3661 && in <= 3665) out = 2906;
	 	 	 else if (in >= 3666 && in <= 3670) out = 2907;
	 	 	 else if (in >= 3671 && in <= 3675) out = 2908;
	 	 	 else if (in >= 3676 && in <= 3679) out = 2909;
	 	 	 else if (in >= 3680 && in <= 3684) out = 2910;
	 	 	 else if (in >= 3685 && in <= 3689) out = 2911;
	 	 	 else if (in >= 3690 && in <= 3694) out = 2912;
	 	 	 else if (in >= 3695 && in <= 3699) out = 2913;
	 	 	 else if (in >= 3700 && in <= 3704) out = 2914;
	 	 	 else if (in >= 3705 && in <= 3709) out = 2915;
	 	 	 else if (in >= 3710 && in <= 3713) out = 2916;
	 	 	 else if (in >= 3714 && in <= 3718) out = 2917;
	 	 	 else if (in >= 3719 && in <= 3723) out = 2918;
	 	 	 else if (in >= 3724 && in <= 3728) out = 2919;
	 	 	 else if (in >= 3729 && in <= 3733) out = 2920;
	 	 	 else if (in >= 3734 && in <= 3738) out = 2921;
	 	 	 else if (in >= 3739 && in <= 3743) out = 2922;
	 	 	 else if (in >= 3744 && in <= 3748) out = 2923;
	 	 	 else if (in >= 3749 && in <= 3753) out = 2924;
	 	 	 else if (in >= 3754 && in <= 3758) out = 2925;
	 	 	 else if (in >= 3759 && in <= 3762) out = 2926;
	 	 	 else if (in >= 3763 && in <= 3767) out = 2927;
	 	 	 else if (in >= 3768 && in <= 3772) out = 2928;
	 	 	 else if (in >= 3773 && in <= 3777) out = 2929;
	 	 	 else if (in >= 3778 && in <= 3782) out = 2930;
	 	 	 else if (in >= 3783 && in <= 3787) out = 2931;
	 	 	 else if (in >= 3788 && in <= 3792) out = 2932;
	 	 	 else if (in >= 3793 && in <= 3797) out = 2933;
	 	 	 else if (in >= 3798 && in <= 3802) out = 2934;
	 	 	 else if (in >= 3803 && in <= 3807) out = 2935;
	 	 	 else if (in >= 3808 && in <= 3812) out = 2936;
	 	 	 else if (in >= 3813 && in <= 3817) out = 2937;
	 	 	 else if (in >= 3818 && in <= 3821) out = 2938;
	 	 	 else if (in >= 3822 && in <= 3826) out = 2939;
	 	 	 else if (in >= 3827 && in <= 3831) out = 2940;
	 	 	 else if (in >= 3832 && in <= 3836) out = 2941;
	 	 	 else if (in >= 3837 && in <= 3841) out = 2942;
	 	 	 else if (in >= 3842 && in <= 3846) out = 2943;
	 	 	 else if (in >= 3847 && in <= 3851) out = 2944;
	 	 	 else if (in >= 3852 && in <= 3856) out = 2945;
	 	 	 else if (in >= 3857 && in <= 3861) out = 2946;
	 	 	 else if (in >= 3862 && in <= 3866) out = 2947;
	 	 	 else if (in >= 3867 && in <= 3871) out = 2948;
	 	 	 else if (in >= 3872 && in <= 3876) out = 2949;
	 	 	 else if (in >= 3877 && in <= 3881) out = 2950;
	 	 	 else if (in >= 3882 && in <= 3886) out = 2951;
	 	 	 else if (in >= 3887 && in <= 3891) out = 2952;
	 	 	 else if (in >= 3892 && in <= 3896) out = 2953;
	 	 	 else if (in >= 3897 && in <= 3901) out = 2954;
	 	 	 else if (in >= 3902 && in <= 3906) out = 2955;
	 	 	 else if (in >= 3907 && in <= 3911) out = 2956;
	 	 	 else if (in >= 3912 && in <= 3916) out = 2957;
	 	 	 else if (in >= 3917 && in <= 3921) out = 2958;
	 	 	 else if (in >= 3922 && in <= 3926) out = 2959;
	 	 	 else if (in >= 3927 && in <= 3931) out = 2960;
	 	 	 else if (in >= 3932 && in <= 3936) out = 2961;
	 	 	 else if (in >= 3937 && in <= 3941) out = 2962;
	 	 	 else if (in >= 3942 && in <= 3946) out = 2963;
	 	 	 else if (in >= 3947 && in <= 3951) out = 2964;
	 	 	 else if (in >= 3952 && in <= 3956) out = 2965;
	 	 	 else if (in >= 3957 && in <= 3961) out = 2966;
	 	 	 else if (in >= 3962 && in <= 3966) out = 2967;
	 	 	 else if (in >= 3967 && in <= 3971) out = 2968;
	 	 	 else if (in >= 3972 && in <= 3976) out = 2969;
	 	 	 else if (in >= 3977 && in <= 3981) out = 2970;
	 	 	 else if (in >= 3982 && in <= 3986) out = 2971;
	 	 	 else if (in >= 3987 && in <= 3991) out = 2972;
	 	 	 else if (in >= 3992 && in <= 3996) out = 2973;
	 	 	 else if (in >= 3997 && in <= 4001) out = 2974;
	 	 	 else if (in >= 4002 && in <= 4006) out = 2975;
	 	 	 else if (in >= 4007 && in <= 4011) out = 2976;
	 	 	 else if (in >= 4012 && in <= 4016) out = 2977;
	 	 	 else if (in >= 4017 && in <= 4021) out = 2978;
	 	 	 else if (in >= 4022 && in <= 4026) out = 2979;
	 	 	 else if (in >= 4027 && in <= 4031) out = 2980;
	 	 	 else if (in >= 4032 && in <= 4036) out = 2981;
	 	 	 else if (in >= 4037 && in <= 4041) out = 2982;
	 	 	 else if (in >= 4042 && in <= 4046) out = 2983;
	 	 	 else if (in >= 4047 && in <= 4051) out = 2984;
	 	 	 else if (in >= 4052 && in <= 4056) out = 2985;
	 	 	 else if (in >= 4057 && in <= 4062) out = 2986;
	 	 	 else if (in >= 4063 && in <= 4067) out = 2987;
	 	 	 else if (in >= 4068 && in <= 4072) out = 2988;
	 	 	 else if (in >= 4073 && in <= 4077) out = 2989;
	 	 	 else if (in >= 4078 && in <= 4082) out = 2990;
	 	 	 else if (in >= 4083 && in <= 4087) out = 2991;
	 	 	 else if (in >= 4088 && in <= 4092) out = 2992;
	 	 	 else if (in >= 4093 && in <= 4097) out = 2993;
	 	 	 else if (in >= 4098 && in <= 4102) out = 2994;
	 	 	 else if (in >= 4103 && in <= 4107) out = 2995;
	 	 	 else if (in >= 4108 && in <= 4112) out = 2996;
	 	 	 else if (in >= 4113 && in <= 4117) out = 2997;
	 	 	 else if (in >= 4118 && in <= 4123) out = 2998;
	 	 	 else if (in >= 4124 && in <= 4128) out = 2999;
	 	 	 else if (in >= 4129 && in <= 4133) out = 3000;
	 	 	 else if (in >= 4134 && in <= 4138) out = 3001;
	 	 	 else if (in >= 4139 && in <= 4143) out = 3002;
	 	 	 else if (in >= 4144 && in <= 4148) out = 3003;
	 	 	 else if (in >= 4149 && in <= 4153) out = 3004;
	 	 	 else if (in >= 4154 && in <= 4158) out = 3005;
	 	 	 else if (in >= 4159 && in <= 4164) out = 3006;
	 	 	 else if (in >= 4165 && in <= 4169) out = 3007;
	 	 	 else if (in >= 4170 && in <= 4174) out = 3008;
	 	 	 else if (in >= 4175 && in <= 4179) out = 3009;
	 	 	 else if (in >= 4180 && in <= 4184) out = 3010;
	 	 	 else if (in >= 4185 && in <= 4189) out = 3011;
	 	 	 else if (in >= 4190 && in <= 4194) out = 3012;
	 	 	 else if (in >= 4195 && in <= 4199) out = 3013;
	 	 	 else if (in >= 4200 && in <= 4205) out = 3014;
	 	 	 else if (in >= 4206 && in <= 4210) out = 3015;
	 	 	 else if (in >= 4211 && in <= 4215) out = 3016;
	 	 	 else if (in >= 4216 && in <= 4220) out = 3017;
	 	 	 else if (in >= 4221 && in <= 4225) out = 3018;
	 	 	 else if (in >= 4226 && in <= 4230) out = 3019;
	 	 	 else if (in >= 4231 && in <= 4236) out = 3020;
	 	 	 else if (in >= 4237 && in <= 4241) out = 3021;
	 	 	 else if (in >= 4242 && in <= 4246) out = 3022;
	 	 	 else if (in >= 4247 && in <= 4251) out = 3023;
	 	 	 else if (in >= 4252 && in <= 4256) out = 3024;
	 	 	 else if (in >= 4257 && in <= 4261) out = 3025;
	 	 	 else if (in >= 4262 && in <= 4267) out = 3026;
	 	 	 else if (in >= 4268 && in <= 4272) out = 3027;
	 	 	 else if (in >= 4273 && in <= 4277) out = 3028;
	 	 	 else if (in >= 4278 && in <= 4282) out = 3029;
	 	 	 else if (in >= 4283 && in <= 4287) out = 3030;
	 	 	 else if (in >= 4288 && in <= 4293) out = 3031;
	 	 	 else if (in >= 4294 && in <= 4298) out = 3032;
	 	 	 else if (in >= 4299 && in <= 4303) out = 3033;
	 	 	 else if (in >= 4304 && in <= 4308) out = 3034;
	 	 	 else if (in >= 4309 && in <= 4313) out = 3035;
	 	 	 else if (in >= 4314 && in <= 4319) out = 3036;
	 	 	 else if (in >= 4320 && in <= 4324) out = 3037;
	 	 	 else if (in >= 4325 && in <= 4329) out = 3038;
	 	 	 else if (in >= 4330 && in <= 4334) out = 3039;
	 	 	 else if (in >= 4335 && in <= 4340) out = 3040;
	 	 	 else if (in >= 4341 && in <= 4345) out = 3041;
	 	 	 else if (in >= 4346 && in <= 4350) out = 3042;
	 	 	 else if (in >= 4351 && in <= 4355) out = 3043;
	 	 	 else if (in >= 4356 && in <= 4361) out = 3044;
	 	 	 else if (in >= 4362 && in <= 4366) out = 3045;
	 	 	 else if (in >= 4367 && in <= 4371) out = 3046;
	 	 	 else if (in >= 4372 && in <= 4376) out = 3047;
	 	 	 else if (in >= 4377 && in <= 4382) out = 3048;
	 	 	 else if (in >= 4383 && in <= 4387) out = 3049;
	 	 	 else if (in >= 4388 && in <= 4392) out = 3050;
	 	 	 else if (in >= 4393 && in <= 4397) out = 3051;
	 	 	 else if (in >= 4398 && in <= 4403) out = 3052;
	 	 	 else if (in >= 4404 && in <= 4408) out = 3053;
	 	 	 else if (in >= 4409 && in <= 4413) out = 3054;
	 	 	 else if (in >= 4414 && in <= 4418) out = 3055;
	 	 	 else if (in >= 4419 && in <= 4424) out = 3056;
	 	 	 else if (in >= 4425 && in <= 4429) out = 3057;
	 	 	 else if (in >= 4430 && in <= 4434) out = 3058;
	 	 	 else if (in >= 4435 && in <= 4440) out = 3059;
	 	 	 else if (in >= 4441 && in <= 4445) out = 3060;
	 	 	 else if (in >= 4446 && in <= 4450) out = 3061;
	 	 	 else if (in >= 4451 && in <= 4456) out = 3062;
	 	 	 else if (in >= 4457 && in <= 4461) out = 3063;
	 	 	 else if (in >= 4462 && in <= 4466) out = 3064;
	 	 	 else if (in >= 4467 && in <= 4471) out = 3065;
	 	 	 else if (in >= 4472 && in <= 4477) out = 3066;
	 	 	 else if (in >= 4478 && in <= 4482) out = 3067;
	 	 	 else if (in >= 4483 && in <= 4487) out = 3068;
	 	 	 else if (in >= 4488 && in <= 4493) out = 3069;
	 	 	 else if (in >= 4494 && in <= 4498) out = 3070;
	 	 	 else if (in >= 4499 && in <= 4503) out = 3071;
	 	 	 else if (in >= 4504 && in <= 4509) out = 3072;
	 	 	 else if (in >= 4510 && in <= 4514) out = 3073;
	 	 	 else if (in >= 4515 && in <= 4519) out = 3074;
	 	 	 else if (in >= 4520 && in <= 4525) out = 3075;
	 	 	 else if (in >= 4526 && in <= 4530) out = 3076;
	 	 	 else if (in >= 4531 && in <= 4536) out = 3077;
	 	 	 else if (in >= 4537 && in <= 4541) out = 3078;
	 	 	 else if (in >= 4542 && in <= 4546) out = 3079;
	 	 	 else if (in >= 4547 && in <= 4552) out = 3080;
	 	 	 else if (in >= 4553 && in <= 4557) out = 3081;
	 	 	 else if (in >= 4558 && in <= 4562) out = 3082;
	 	 	 else if (in >= 4563 && in <= 4568) out = 3083;
	 	 	 else if (in >= 4569 && in <= 4573) out = 3084;
	 	 	 else if (in >= 4574 && in <= 4578) out = 3085;
	 	 	 else if (in >= 4579 && in <= 4584) out = 3086;
	 	 	 else if (in >= 4585 && in <= 4589) out = 3087;
	 	 	 else if (in >= 4590 && in <= 4595) out = 3088;
	 	 	 else if (in >= 4596 && in <= 4600) out = 3089;
	 	 	 else if (in >= 4601 && in <= 4605) out = 3090;
	 	 	 else if (in >= 4606 && in <= 4611) out = 3091;
	 	 	 else if (in >= 4612 && in <= 4616) out = 3092;
	 	 	 else if (in >= 4617 && in <= 4622) out = 3093;
	 	 	 else if (in >= 4623 && in <= 4627) out = 3094;
	 	 	 else if (in >= 4628 && in <= 4633) out = 3095;
	 	 	 else if (in >= 4634 && in <= 4638) out = 3096;
	 	 	 else if (in >= 4639 && in <= 4643) out = 3097;
	 	 	 else if (in >= 4644 && in <= 4649) out = 3098;
	 	 	 else if (in >= 4650 && in <= 4654) out = 3099;
	 	 	 else if (in >= 4655 && in <= 4660) out = 3100;
	 	 	 else if (in >= 4661 && in <= 4665) out = 3101;
	 	 	 else if (in >= 4666 && in <= 4671) out = 3102;
	 	 	 else if (in >= 4672 && in <= 4676) out = 3103;
	 	 	 else if (in >= 4677 && in <= 4681) out = 3104;
	 	 	 else if (in >= 4682 && in <= 4687) out = 3105;
	 	 	 else if (in >= 4688 && in <= 4692) out = 3106;
	 	 	 else if (in >= 4693 && in <= 4698) out = 3107;
	 	 	 else if (in >= 4699 && in <= 4703) out = 3108;
	 	 	 else if (in >= 4704 && in <= 4709) out = 3109;
	 	 	 else if (in >= 4710 && in <= 4714) out = 3110;
	 	 	 else if (in >= 4715 && in <= 4720) out = 3111;
	 	 	 else if (in >= 4721 && in <= 4725) out = 3112;
	 	 	 else if (in >= 4726 && in <= 4731) out = 3113;
	 	 	 else if (in >= 4732 && in <= 4736) out = 3114;
	 	 	 else if (in >= 4737 && in <= 4742) out = 3115;
	 	 	 else if (in >= 4743 && in <= 4747) out = 3116;
	 	 	 else if (in >= 4748 && in <= 4753) out = 3117;
	 	 	 else if (in >= 4754 && in <= 4758) out = 3118;
	 	 	 else if (in >= 4759 && in <= 4764) out = 3119;
	 	 	 else if (in >= 4765 && in <= 4769) out = 3120;
	 	 	 else if (in >= 4770 && in <= 4775) out = 3121;
	 	 	 else if (in >= 4776 && in <= 4780) out = 3122;
	 	 	 else if (in >= 4781 && in <= 4786) out = 3123;
	 	 	 else if (in >= 4787 && in <= 4791) out = 3124;
	 	 	 else if (in >= 4792 && in <= 4797) out = 3125;
	 	 	 else if (in >= 4798 && in <= 4802) out = 3126;
	 	 	 else if (in >= 4803 && in <= 4808) out = 3127;
	 	 	 else if (in >= 4809 && in <= 4814) out = 3128;
	 	 	 else if (in >= 4815 && in <= 4819) out = 3129;
	 	 	 else if (in >= 4820 && in <= 4825) out = 3130;
	 	 	 else if (in >= 4826 && in <= 4830) out = 3131;
	 	 	 else if (in >= 4831 && in <= 4836) out = 3132;
	 	 	 else if (in >= 4837 && in <= 4841) out = 3133;
	 	 	 else if (in >= 4842 && in <= 4847) out = 3134;
	 	 	 else if (in >= 4848 && in <= 4852) out = 3135;
	 	 	 else if (in >= 4853 && in <= 4858) out = 3136;
	 	 	 else if (in >= 4859 && in <= 4864) out = 3137;
	 	 	 else if (in >= 4865 && in <= 4869) out = 3138;
	 	 	 else if (in >= 4870 && in <= 4875) out = 3139;
	 	 	 else if (in >= 4876 && in <= 4880) out = 3140;
	 	 	 else if (in >= 4881 && in <= 4886) out = 3141;
	 	 	 else if (in >= 4887 && in <= 4892) out = 3142;
	 	 	 else if (in >= 4893 && in <= 4897) out = 3143;
	 	 	 else if (in >= 4898 && in <= 4903) out = 3144;
	 	 	 else if (in >= 4904 && in <= 4908) out = 3145;
	 	 	 else if (in >= 4909 && in <= 4914) out = 3146;
	 	 	 else if (in >= 4915 && in <= 4920) out = 3147;
	 	 	 else if (in >= 4921 && in <= 4925) out = 3148;
	 	 	 else if (in >= 4926 && in <= 4931) out = 3149;
	 	 	 else if (in >= 4932 && in <= 4937) out = 3150;
	 	 	 else if (in >= 4938 && in <= 4942) out = 3151;
	 	 	 else if (in >= 4943 && in <= 4948) out = 3152;
	 	 	 else if (in >= 4949 && in <= 4954) out = 3153;
	 	 	 else if (in >= 4955 && in <= 4959) out = 3154;
	 	 	 else if (in >= 4960 && in <= 4965) out = 3155;
	 	 	 else if (in >= 4966 && in <= 4971) out = 3156;
	 	 	 else if (in >= 4972 && in <= 4976) out = 3157;
	 	 	 else if (in >= 4977 && in <= 4982) out = 3158;
	 	 	 else if (in >= 4983 && in <= 4988) out = 3159;
	 	 	 else if (in >= 4989 && in <= 4993) out = 3160;
	 	 	 else if (in >= 4994 && in <= 4999) out = 3161;
	 	 	 else if (in >= 5000 && in <= 5005) out = 3162;
	 	 	 else if (in >= 5006 && in <= 5010) out = 3163;
	 	 	 else if (in >= 5011 && in <= 5016) out = 3164;
	 	 	 else if (in >= 5017 && in <= 5022) out = 3165;
	 	 	 else if (in >= 5023 && in <= 5027) out = 3166;
	 	 	 else if (in >= 5028 && in <= 5033) out = 3167;
	 	 	 else if (in >= 5034 && in <= 5039) out = 3168;
	 	 	 else if (in >= 5040 && in <= 5045) out = 3169;
	 	 	 else if (in >= 5046 && in <= 5050) out = 3170;
	 	 	 else if (in >= 5051 && in <= 5056) out = 3171;
	 	 	 else if (in >= 5057 && in <= 5062) out = 3172;
	 	 	 else if (in >= 5063 && in <= 5067) out = 3173;
	 	 	 else if (in >= 5068 && in <= 5073) out = 3174;
	 	 	 else if (in >= 5074 && in <= 5079) out = 3175;
	 	 	 else if (in >= 5080 && in <= 5085) out = 3176;
	 	 	 else if (in >= 5086 && in <= 5090) out = 3177;
	 	 	 else if (in >= 5091 && in <= 5096) out = 3178;
	 	 	 else if (in >= 5097 && in <= 5102) out = 3179;
	 	 	 else if (in >= 5103 && in <= 5108) out = 3180;
	 	 	 else if (in >= 5109 && in <= 5113) out = 3181;
	 	 	 else if (in >= 5114 && in <= 5119) out = 3182;
	 	 	 else if (in >= 5120 && in <= 5125) out = 3183;
	 	 	 else if (in >= 5126 && in <= 5131) out = 3184;
	 	 	 else if (in >= 5132 && in <= 5137) out = 3185;
	 	 	 else if (in >= 5138 && in <= 5142) out = 3186;
	 	 	 else if (in >= 5143 && in <= 5148) out = 3187;
	 	 	 else if (in >= 5149 && in <= 5154) out = 3188;
	 	 	 else if (in >= 5155 && in <= 5160) out = 3189;
	 	 	 else if (in >= 5161 && in <= 5166) out = 3190;
	 	 	 else if (in >= 5167 && in <= 5171) out = 3191;
	 	 	 else if (in >= 5172 && in <= 5177) out = 3192;
	 	 	 else if (in >= 5178 && in <= 5183) out = 3193;
	 	 	 else if (in >= 5184 && in <= 5189) out = 3194;
	 	 	 else if (in >= 5190 && in <= 5195) out = 3195;
	 	 	 else if (in >= 5196 && in <= 5201) out = 3196;
	 	 	 else if (in >= 5202 && in <= 5206) out = 3197;
	 	 	 else if (in >= 5207 && in <= 5212) out = 3198;
	 	 	 else if (in >= 5213 && in <= 5218) out = 3199;
	 	 	 else if (in >= 5219 && in <= 5224) out = 3200;
	 	 	 else if (in >= 5225 && in <= 5230) out = 3201;
	 	 	 else if (in >= 5231 && in <= 5236) out = 3202;
	 	 	 else if (in >= 5237 && in <= 5242) out = 3203;
	 	 	 else if (in >= 5243 && in <= 5247) out = 3204;
	 	 	 else if (in >= 5248 && in <= 5253) out = 3205;
	 	 	 else if (in >= 5254 && in <= 5259) out = 3206;
	 	 	 else if (in >= 5260 && in <= 5265) out = 3207;
	 	 	 else if (in >= 5266 && in <= 5271) out = 3208;
	 	 	 else if (in >= 5272 && in <= 5277) out = 3209;
	 	 	 else if (in >= 5278 && in <= 5283) out = 3210;
	 	 	 else if (in >= 5284 && in <= 5289) out = 3211;
	 	 	 else if (in >= 5290 && in <= 5295) out = 3212;
	 	 	 else if (in >= 5296 && in <= 5301) out = 3213;
	 	 	 else if (in >= 5302 && in <= 5307) out = 3214;
	 	 	 else if (in >= 5308 && in <= 5312) out = 3215;
	 	 	 else if (in >= 5313 && in <= 5318) out = 3216;
	 	 	 else if (in >= 5319 && in <= 5324) out = 3217;
	 	 	 else if (in >= 5325 && in <= 5330) out = 3218;
	 	 	 else if (in >= 5331 && in <= 5336) out = 3219;
	 	 	 else if (in >= 5337 && in <= 5342) out = 3220;
	 	 	 else if (in >= 5343 && in <= 5348) out = 3221;
	 	 	 else if (in >= 5349 && in <= 5354) out = 3222;
	 	 	 else if (in >= 5355 && in <= 5360) out = 3223;
	 	 	 else if (in >= 5361 && in <= 5366) out = 3224;
	 	 	 else if (in >= 5367 && in <= 5372) out = 3225;
	 	 	 else if (in >= 5373 && in <= 5378) out = 3226;
	 	 	 else if (in >= 5379 && in <= 5384) out = 3227;
	 	 	 else if (in >= 5385 && in <= 5390) out = 3228;
	 	 	 else if (in >= 5391 && in <= 5396) out = 3229;
	 	 	 else if (in >= 5397 && in <= 5402) out = 3230;
	 	 	 else if (in >= 5403 && in <= 5408) out = 3231;
	 	 	 else if (in >= 5409 && in <= 5414) out = 3232;
	 	 	 else if (in >= 5415 && in <= 5420) out = 3233;
	 	 	 else if (in >= 5421 && in <= 5426) out = 3234;
	 	 	 else if (in >= 5427 && in <= 5432) out = 3235;
	 	 	 else if (in >= 5433 && in <= 5438) out = 3236;
	 	 	 else if (in >= 5439 && in <= 5444) out = 3237;
	 	 	 else if (in >= 5445 && in <= 5450) out = 3238;
	 	 	 else if (in >= 5451 && in <= 5456) out = 3239;
	 	 	 else if (in >= 5457 && in <= 5462) out = 3240;
	 	 	 else if (in >= 5463 && in <= 5468) out = 3241;
	 	 	 else if (in >= 5469 && in <= 5474) out = 3242;
	 	 	 else if (in >= 5475 && in <= 5481) out = 3243;
	 	 	 else if (in >= 5482 && in <= 5487) out = 3244;
	 	 	 else if (in >= 5488 && in <= 5493) out = 3245;
	 	 	 else if (in >= 5494 && in <= 5499) out = 3246;
	 	 	 else if (in >= 5500 && in <= 5505) out = 3247;
	 	 	 else if (in >= 5506 && in <= 5511) out = 3248;
	 	 	 else if (in >= 5512 && in <= 5517) out = 3249;
	 	 	 else if (in >= 5518 && in <= 5523) out = 3250;
	 	 	 else if (in >= 5524 && in <= 5529) out = 3251;
	 	 	 else if (in >= 5530 && in <= 5535) out = 3252;
	 	 	 else if (in >= 5536 && in <= 5542) out = 3253;
	 	 	 else if (in >= 5543 && in <= 5548) out = 3254;
	 	 	 else if (in >= 5549 && in <= 5554) out = 3255;
	 	 	 else if (in >= 5555 && in <= 5560) out = 3256;
	 	 	 else if (in >= 5561 && in <= 5566) out = 3257;
	 	 	 else if (in >= 5567 && in <= 5572) out = 3258;
	 	 	 else if (in >= 5573 && in <= 5578) out = 3259;
	 	 	 else if (in >= 5579 && in <= 5585) out = 3260;
	 	 	 else if (in >= 5586 && in <= 5591) out = 3261;
	 	 	 else if (in >= 5592 && in <= 5597) out = 3262;
	 	 	 else if (in >= 5598 && in <= 5603) out = 3263;
	 	 	 else if (in >= 5604 && in <= 5609) out = 3264;
	 	 	 else if (in >= 5610 && in <= 5616) out = 3265;
	 	 	 else if (in >= 5617 && in <= 5622) out = 3266;
	 	 	 else if (in >= 5623 && in <= 5628) out = 3267;
	 	 	 else if (in >= 5629 && in <= 5634) out = 3268;
	 	 	 else if (in >= 5635 && in <= 5640) out = 3269;
	 	 	 else if (in >= 5641 && in <= 5647) out = 3270;
	 	 	 else if (in >= 5648 && in <= 5653) out = 3271;
	 	 	 else if (in >= 5654 && in <= 5659) out = 3272;
	 	 	 else if (in >= 5660 && in <= 5665) out = 3273;
	 	 	 else if (in >= 5666 && in <= 5672) out = 3274;
	 	 	 else if (in >= 5673 && in <= 5678) out = 3275;
	 	 	 else if (in >= 5679 && in <= 5684) out = 3276;
	 	 	 else if (in >= 5685 && in <= 5690) out = 3277;
	 	 	 else if (in >= 5691 && in <= 5697) out = 3278;
	 	 	 else if (in >= 5698 && in <= 5703) out = 3279;
	 	 	 else if (in >= 5704 && in <= 5709) out = 3280;
	 	 	 else if (in >= 5710 && in <= 5715) out = 3281;
	 	 	 else if (in >= 5716 && in <= 5722) out = 3282;
	 	 	 else if (in >= 5723 && in <= 5728) out = 3283;
	 	 	 else if (in >= 5729 && in <= 5734) out = 3284;
	 	 	 else if (in >= 5735 && in <= 5741) out = 3285;
	 	 	 else if (in >= 5742 && in <= 5747) out = 3286;
	 	 	 else if (in >= 5748 && in <= 5753) out = 3287;
	 	 	 else if (in >= 5754 && in <= 5760) out = 3288;
	 	 	 else if (in >= 5761 && in <= 5766) out = 3289;
	 	 	 else if (in >= 5767 && in <= 5772) out = 3290;
	 	 	 else if (in >= 5773 && in <= 5779) out = 3291;
	 	 	 else if (in >= 5780 && in <= 5785) out = 3292;
	 	 	 else if (in >= 5786 && in <= 5791) out = 3293;
	 	 	 else if (in >= 5792 && in <= 5798) out = 3294;
	 	 	 else if (in >= 5799 && in <= 5804) out = 3295;
	 	 	 else if (in >= 5805 && in <= 5810) out = 3296;
	 	 	 else if (in >= 5811 && in <= 5817) out = 3297;
	 	 	 else if (in >= 5818 && in <= 5823) out = 3298;
	 	 	 else if (in >= 5824 && in <= 5829) out = 3299;
	 	 	 else if (in >= 5830 && in <= 5836) out = 3300;
	 	 	 else if (in >= 5837 && in <= 5842) out = 3301;
	 	 	 else if (in >= 5843 && in <= 5849) out = 3302;
	 	 	 else if (in >= 5850 && in <= 5855) out = 3303;
	 	 	 else if (in >= 5856 && in <= 5862) out = 3304;
	 	 	 else if (in >= 5863 && in <= 5868) out = 3305;
	 	 	 else if (in >= 5869 && in <= 5874) out = 3306;
	 	 	 else if (in >= 5875 && in <= 5881) out = 3307;
	 	 	 else if (in >= 5882 && in <= 5887) out = 3308;
	 	 	 else if (in >= 5888 && in <= 5894) out = 3309;
	 	 	 else if (in >= 5895 && in <= 5900) out = 3310;
	 	 	 else if (in >= 5901 && in <= 5907) out = 3311;
	 	 	 else if (in >= 5908 && in <= 5913) out = 3312;
	 	 	 else if (in >= 5914 && in <= 5920) out = 3313;
	 	 	 else if (in >= 5921 && in <= 5926) out = 3314;
	 	 	 else if (in >= 5927 && in <= 5933) out = 3315;
	 	 	 else if (in >= 5934 && in <= 5939) out = 3316;
	 	 	 else if (in >= 5940 && in <= 5946) out = 3317;
	 	 	 else if (in >= 5947 && in <= 5952) out = 3318;
	 	 	 else if (in >= 5953 && in <= 5959) out = 3319;
	 	 	 else if (in >= 5960 && in <= 5965) out = 3320;
	 	 	 else if (in >= 5966 && in <= 5972) out = 3321;
	 	 	 else if (in >= 5973 && in <= 5978) out = 3322;
	 	 	 else if (in >= 5979 && in <= 5985) out = 3323;
	 	 	 else if (in >= 5986 && in <= 5991) out = 3324;
	 	 	 else if (in >= 5992 && in <= 5998) out = 3325;
	 	 	 else if (in >= 5999 && in <= 6004) out = 3326;
	 	 	 else if (in >= 6005 && in <= 6011) out = 3327;
	 	 	 else if (in >= 6012 && in <= 6018) out = 3328;
	 	 	 else if (in >= 6019 && in <= 6024) out = 3329;
	 	 	 else if (in >= 6025 && in <= 6031) out = 3330;
	 	 	 else if (in >= 6032 && in <= 6037) out = 3331;
	 	 	 else if (in >= 6038 && in <= 6044) out = 3332;
	 	 	 else if (in >= 6045 && in <= 6050) out = 3333;
	 	 	 else if (in >= 6051 && in <= 6057) out = 3334;
	 	 	 else if (in >= 6058 && in <= 6064) out = 3335;
	 	 	 else if (in >= 6065 && in <= 6070) out = 3336;
	 	 	 else if (in >= 6071 && in <= 6077) out = 3337;
	 	 	 else if (in >= 6078 && in <= 6084) out = 3338;
	 	 	 else if (in >= 6085 && in <= 6090) out = 3339;
	 	 	 else if (in >= 6091 && in <= 6097) out = 3340;
	 	 	 else if (in >= 6098 && in <= 6104) out = 3341;
	 	 	 else if (in >= 6105 && in <= 6110) out = 3342;
	 	 	 else if (in >= 6111 && in <= 6117) out = 3343;
	 	 	 else if (in >= 6118 && in <= 6124) out = 3344;
	 	 	 else if (in >= 6125 && in <= 6130) out = 3345;
	 	 	 else if (in >= 6131 && in <= 6137) out = 3346;
	 	 	 else if (in >= 6138 && in <= 6144) out = 3347;
	 	 	 else if (in >= 6145 && in <= 6150) out = 3348;
	 	 	 else if (in >= 6151 && in <= 6157) out = 3349;
	 	 	 else if (in >= 6158 && in <= 6164) out = 3350;
	 	 	 else if (in >= 6165 && in <= 6171) out = 3351;
	 	 	 else if (in >= 6172 && in <= 6177) out = 3352;
	 	 	 else if (in >= 6178 && in <= 6184) out = 3353;
	 	 	 else if (in >= 6185 && in <= 6191) out = 3354;
	 	 	 else if (in >= 6192 && in <= 6198) out = 3355;
	 	 	 else if (in >= 6199 && in <= 6204) out = 3356;
	 	 	 else if (in >= 6205 && in <= 6211) out = 3357;
	 	 	 else if (in >= 6212 && in <= 6218) out = 3358;
	 	 	 else if (in >= 6219 && in <= 6225) out = 3359;
	 	 	 else if (in >= 6226 && in <= 6232) out = 3360;
	 	 	 else if (in >= 6233 && in <= 6238) out = 3361;
	 	 	 else if (in >= 6239 && in <= 6245) out = 3362;
	 	 	 else if (in >= 6246 && in <= 6252) out = 3363;
	 	 	 else if (in >= 6253 && in <= 6259) out = 3364;
	 	 	 else if (in >= 6260 && in <= 6266) out = 3365;
	 	 	 else if (in >= 6267 && in <= 6272) out = 3366;
	 	 	 else if (in >= 6273 && in <= 6279) out = 3367;
	 	 	 else if (in >= 6280 && in <= 6286) out = 3368;
	 	 	 else if (in >= 6287 && in <= 6293) out = 3369;
	 	 	 else if (in >= 6294 && in <= 6300) out = 3370;
	 	 	 else if (in >= 6301 && in <= 6307) out = 3371;
	 	 	 else if (in >= 6308 && in <= 6314) out = 3372;
	 	 	 else if (in >= 6315 && in <= 6321) out = 3373;
	 	 	 else if (in >= 6322 && in <= 6327) out = 3374;
	 	 	 else if (in >= 6328 && in <= 6334) out = 3375;
	 	 	 else if (in >= 6335 && in <= 6341) out = 3376;
	 	 	 else if (in >= 6342 && in <= 6348) out = 3377;
	 	 	 else if (in >= 6349 && in <= 6355) out = 3378;
	 	 	 else if (in >= 6356 && in <= 6362) out = 3379;
	 	 	 else if (in >= 6363 && in <= 6369) out = 3380;
	 	 	 else if (in >= 6370 && in <= 6376) out = 3381;
	 	 	 else if (in >= 6377 && in <= 6383) out = 3382;
	 	 	 else if (in >= 6384 && in <= 6390) out = 3383;
	 	 	 else if (in >= 6391 && in <= 6397) out = 3384;
	 	 	 else if (in >= 6398 && in <= 6404) out = 3385;
	 	 	 else if (in >= 6405 && in <= 6411) out = 3386;
	 	 	 else if (in >= 6412 && in <= 6418) out = 3387;
	 	 	 else if (in >= 6419 && in <= 6425) out = 3388;
	 	 	 else if (in >= 6426 && in <= 6432) out = 3389;
	 	 	 else if (in >= 6433 && in <= 6439) out = 3390;
	 	 	 else if (in >= 6440 && in <= 6446) out = 3391;
	 	 	 else if (in >= 6447 && in <= 6453) out = 3392;
	 	 	 else if (in >= 6454 && in <= 6460) out = 3393;
	 	 	 else if (in >= 6461 && in <= 6467) out = 3394;
	 	 	 else if (in >= 6468 && in <= 6474) out = 3395;
	 	 	 else if (in >= 6475 && in <= 6481) out = 3396;
	 	 	 else if (in >= 6482 && in <= 6488) out = 3397;
	 	 	 else if (in >= 6489 && in <= 6495) out = 3398;
	 	 	 else if (in >= 6496 && in <= 6502) out = 3399;
	 	 	 else if (in >= 6503 && in <= 6509) out = 3400;
	 	 	 else if (in >= 6510 && in <= 6517) out = 3401;
	 	 	 else if (in >= 6518 && in <= 6524) out = 3402;
	 	 	 else if (in >= 6525 && in <= 6531) out = 3403;
	 	 	 else if (in >= 6532 && in <= 6538) out = 3404;
	 	 	 else if (in >= 6539 && in <= 6545) out = 3405;
	 	 	 else if (in >= 6546 && in <= 6552) out = 3406;
	 	 	 else if (in >= 6553 && in <= 6559) out = 3407;
	 	 	 else if (in >= 6560 && in <= 6567) out = 3408;
	 	 	 else if (in >= 6568 && in <= 6574) out = 3409;
	 	 	 else if (in >= 6575 && in <= 6581) out = 3410;
	 	 	 else if (in >= 6582 && in <= 6588) out = 3411;
	 	 	 else if (in >= 6589 && in <= 6595) out = 3412;
	 	 	 else if (in >= 6596 && in <= 6603) out = 3413;
	 	 	 else if (in >= 6604 && in <= 6610) out = 3414;
	 	 	 else if (in >= 6611 && in <= 6617) out = 3415;
	 	 	 else if (in >= 6618 && in <= 6624) out = 3416;
	 	 	 else if (in >= 6625 && in <= 6631) out = 3417;
	 	 	 else if (in >= 6632 && in <= 6639) out = 3418;
	 	 	 else if (in >= 6640 && in <= 6646) out = 3419;
	 	 	 else if (in >= 6647 && in <= 6653) out = 3420;
	 	 	 else if (in >= 6654 && in <= 6661) out = 3421;
	 	 	 else if (in >= 6662 && in <= 6668) out = 3422;
	 	 	 else if (in >= 6669 && in <= 6675) out = 3423;
	 	 	 else if (in >= 6676 && in <= 6682) out = 3424;
	 	 	 else if (in >= 6683 && in <= 6690) out = 3425;
	 	 	 else if (in >= 6691 && in <= 6697) out = 3426;
	 	 	 else if (in >= 6698 && in <= 6704) out = 3427;
	 	 	 else if (in >= 6705 && in <= 6712) out = 3428;
	 	 	 else if (in >= 6713 && in <= 6719) out = 3429;
	 	 	 else if (in >= 6720 && in <= 6726) out = 3430;
	 	 	 else if (in >= 6727 && in <= 6734) out = 3431;
	 	 	 else if (in >= 6735 && in <= 6741) out = 3432;
	 	 	 else if (in >= 6742 && in <= 6749) out = 3433;
	 	 	 else if (in >= 6750 && in <= 6756) out = 3434;
	 	 	 else if (in >= 6757 && in <= 6763) out = 3435;
	 	 	 else if (in >= 6764 && in <= 6771) out = 3436;
	 	 	 else if (in >= 6772 && in <= 6778) out = 3437;
	 	 	 else if (in >= 6779 && in <= 6786) out = 3438;
	 	 	 else if (in >= 6787 && in <= 6793) out = 3439;
	 	 	 else if (in >= 6794 && in <= 6801) out = 3440;
	 	 	 else if (in >= 6802 && in <= 6808) out = 3441;
	 	 	 else if (in >= 6809 && in <= 6815) out = 3442;
	 	 	 else if (in >= 6816 && in <= 6823) out = 3443;
	 	 	 else if (in >= 6824 && in <= 6830) out = 3444;
	 	 	 else if (in >= 6831 && in <= 6838) out = 3445;
	 	 	 else if (in >= 6839 && in <= 6845) out = 3446;
	 	 	 else if (in >= 6846 && in <= 6853) out = 3447;
	 	 	 else if (in >= 6854 && in <= 6860) out = 3448;
	 	 	 else if (in >= 6861 && in <= 6868) out = 3449;
	 	 	 else if (in >= 6869 && in <= 6876) out = 3450;
	 	 	 else if (in >= 6877 && in <= 6883) out = 3451;
	 	 	 else if (in >= 6884 && in <= 6891) out = 3452;
	 	 	 else if (in >= 6892 && in <= 6898) out = 3453;
	 	 	 else if (in >= 6899 && in <= 6906) out = 3454;
	 	 	 else if (in >= 6907 && in <= 6913) out = 3455;
	 	 	 else if (in >= 6914 && in <= 6921) out = 3456;
	 	 	 else if (in >= 6922 && in <= 6929) out = 3457;
	 	 	 else if (in >= 6930 && in <= 6936) out = 3458;
	 	 	 else if (in >= 6937 && in <= 6944) out = 3459;
	 	 	 else if (in >= 6945 && in <= 6951) out = 3460;
	 	 	 else if (in >= 6952 && in <= 6959) out = 3461;
	 	 	 else if (in >= 6960 && in <= 6967) out = 3462;
	 	 	 else if (in >= 6968 && in <= 6974) out = 3463;
	 	 	 else if (in >= 6975 && in <= 6982) out = 3464;
	 	 	 else if (in >= 6983 && in <= 6990) out = 3465;
	 	 	 else if (in >= 6991 && in <= 6998) out = 3466;
	 	 	 else if (in >= 6999 && in <= 7005) out = 3467;
	 	 	 else if (in >= 7006 && in <= 7013) out = 3468;
	 	 	 else if (in >= 7014 && in <= 7021) out = 3469;
	 	 	 else if (in >= 7022 && in <= 7028) out = 3470;
	 	 	 else if (in >= 7029 && in <= 7036) out = 3471;
	 	 	 else if (in >= 7037 && in <= 7044) out = 3472;
	 	 	 else if (in >= 7045 && in <= 7052) out = 3473;
	 	 	 else if (in >= 7053 && in <= 7059) out = 3474;
	 	 	 else if (in >= 7060 && in <= 7067) out = 3475;
	 	 	 else if (in >= 7068 && in <= 7075) out = 3476;
	 	 	 else if (in >= 7076 && in <= 7083) out = 3477;
	 	 	 else if (in >= 7084 && in <= 7091) out = 3478;
	 	 	 else if (in >= 7092 && in <= 7099) out = 3479;
	 	 	 else if (in >= 7100 && in <= 7106) out = 3480;
	 	 	 else if (in >= 7107 && in <= 7114) out = 3481;
	 	 	 else if (in >= 7115 && in <= 7122) out = 3482;
	 	 	 else if (in >= 7123 && in <= 7130) out = 3483;
	 	 	 else if (in >= 7131 && in <= 7138) out = 3484;
	 	 	 else if (in >= 7139 && in <= 7146) out = 3485;
	 	 	 else if (in >= 7147 && in <= 7154) out = 3486;
	 	 	 else if (in >= 7155 && in <= 7162) out = 3487;
	 	 	 else if (in >= 7163 && in <= 7170) out = 3488;
	 	 	 else if (in >= 7171 && in <= 7177) out = 3489;
	 	 	 else if (in >= 7178 && in <= 7185) out = 3490;
	 	 	 else if (in >= 7186 && in <= 7193) out = 3491;
	 	 	 else if (in >= 7194 && in <= 7201) out = 3492;
	 	 	 else if (in >= 7202 && in <= 7209) out = 3493;
	 	 	 else if (in >= 7210 && in <= 7217) out = 3494;
	 	 	 else if (in >= 7218 && in <= 7225) out = 3495;
	 	 	 else if (in >= 7226 && in <= 7233) out = 3496;
	 	 	 else if (in >= 7234 && in <= 7241) out = 3497;
	 	 	 else if (in >= 7242 && in <= 7249) out = 3498;
	 	 	 else if (in >= 7250 && in <= 7257) out = 3499;
	 	 	 else if (in >= 7258 && in <= 7265) out = 3500;
	 	 	 else if (in >= 7266 && in <= 7274) out = 3501;
	 	 	 else if (in >= 7275 && in <= 7282) out = 3502;
	 	 	 else if (in >= 7283 && in <= 7290) out = 3503;
	 	 	 else if (in >= 7291 && in <= 7298) out = 3504;
	 	 	 else if (in >= 7299 && in <= 7306) out = 3505;
	 	 	 else if (in >= 7307 && in <= 7314) out = 3506;
	 	 	 else if (in >= 7315 && in <= 7322) out = 3507;
	 	 	 else if (in >= 7323 && in <= 7330) out = 3508;
	 	 	 else if (in >= 7331 && in <= 7339) out = 3509;
	 	 	 else if (in >= 7340 && in <= 7347) out = 3510;
	 	 	 else if (in >= 7348 && in <= 7355) out = 3511;
	 	 	 else if (in >= 7356 && in <= 7363) out = 3512;
	 	 	 else if (in >= 7364 && in <= 7371) out = 3513;
	 	 	 else if (in >= 7372 && in <= 7380) out = 3514;
	 	 	 else if (in >= 7381 && in <= 7388) out = 3515;
	 	 	 else if (in >= 7389 && in <= 7396) out = 3516;
	 	 	 else if (in >= 7397 && in <= 7404) out = 3517;
	 	 	 else if (in >= 7405 && in <= 7413) out = 3518;
	 	 	 else if (in >= 7414 && in <= 7421) out = 3519;
	 	 	 else if (in >= 7422 && in <= 7429) out = 3520;
	 	 	 else if (in >= 7430 && in <= 7437) out = 3521;
	 	 	 else if (in >= 7438 && in <= 7446) out = 3522;
	 	 	 else if (in >= 7447 && in <= 7454) out = 3523;
	 	 	 else if (in >= 7455 && in <= 7462) out = 3524;
	 	 	 else if (in >= 7463 && in <= 7471) out = 3525;
	 	 	 else if (in >= 7472 && in <= 7479) out = 3526;
	 	 	 else if (in >= 7480 && in <= 7488) out = 3527;
	 	 	 else if (in >= 7489 && in <= 7496) out = 3528;
	 	 	 else if (in >= 7497 && in <= 7504) out = 3529;
	 	 	 else if (in >= 7505 && in <= 7513) out = 3530;
	 	 	 else if (in >= 7514 && in <= 7521) out = 3531;
	 	 	 else if (in >= 7522 && in <= 7530) out = 3532;
	 	 	 else if (in >= 7531 && in <= 7538) out = 3533;
	 	 	 else if (in >= 7539 && in <= 7547) out = 3534;
	 	 	 else if (in >= 7548 && in <= 7555) out = 3535;
	 	 	 else if (in >= 7556 && in <= 7563) out = 3536;
	 	 	 else if (in >= 7564 && in <= 7572) out = 3537;
	 	 	 else if (in >= 7573 && in <= 7581) out = 3538;
	 	 	 else if (in >= 7582 && in <= 7589) out = 3539;
	 	 	 else if (in >= 7590 && in <= 7598) out = 3540;
	 	 	 else if (in >= 7599 && in <= 7606) out = 3541;
	 	 	 else if (in >= 7607 && in <= 7615) out = 3542;
	 	 	 else if (in >= 7616 && in <= 7623) out = 3543;
	 	 	 else if (in >= 7624 && in <= 7632) out = 3544;
	 	 	 else if (in >= 7633 && in <= 7640) out = 3545;
	 	 	 else if (in >= 7641 && in <= 7649) out = 3546;
	 	 	 else if (in >= 7650 && in <= 7658) out = 3547;
	 	 	 else if (in >= 7659 && in <= 7666) out = 3548;
	 	 	 else if (in >= 7667 && in <= 7675) out = 3549;
	 	 	 else if (in >= 7676 && in <= 7684) out = 3550;
	 	 	 else if (in >= 7685 && in <= 7692) out = 3551;
	 	 	 else if (in >= 7693 && in <= 7701) out = 3552;
	 	 	 else if (in >= 7702 && in <= 7710) out = 3553;
	 	 	 else if (in >= 7711 && in <= 7719) out = 3554;
	 	 	 else if (in >= 7720 && in <= 7727) out = 3555;
	 	 	 else if (in >= 7728 && in <= 7736) out = 3556;
	 	 	 else if (in >= 7737 && in <= 7745) out = 3557;
	 	 	 else if (in >= 7746 && in <= 7754) out = 3558;
	 	 	 else if (in >= 7755 && in <= 7762) out = 3559;
	 	 	 else if (in >= 7763 && in <= 7771) out = 3560;
	 	 	 else if (in >= 7772 && in <= 7780) out = 3561;
	 	 	 else if (in >= 7781 && in <= 7789) out = 3562;
	 	 	 else if (in >= 7790 && in <= 7798) out = 3563;
	 	 	 else if (in >= 7799 && in <= 7807) out = 3564;
	 	 	 else if (in >= 7808 && in <= 7816) out = 3565;
	 	 	 else if (in >= 7817 && in <= 7824) out = 3566;
	 	 	 else if (in >= 7825 && in <= 7833) out = 3567;
	 	 	 else if (in >= 7834 && in <= 7842) out = 3568;
	 	 	 else if (in >= 7843 && in <= 7851) out = 3569;
	 	 	 else if (in >= 7852 && in <= 7860) out = 3570;
	 	 	 else if (in >= 7861 && in <= 7869) out = 3571;
	 	 	 else if (in >= 7870 && in <= 7878) out = 3572;
	 	 	 else if (in >= 7879 && in <= 7887) out = 3573;
	 	 	 else if (in >= 7888 && in <= 7896) out = 3574;
	 	 	 else if (in >= 7897 && in <= 7905) out = 3575;
	 	 	 else if (in >= 7906 && in <= 7914) out = 3576;
	 	 	 else if (in >= 7915 && in <= 7923) out = 3577;
	 	 	 else if (in >= 7924 && in <= 7932) out = 3578;
	 	 	 else if (in >= 7933 && in <= 7941) out = 3579;
	 	 	 else if (in >= 7942 && in <= 7951) out = 3580;
	 	 	 else if (in >= 7952 && in <= 7960) out = 3581;
	 	 	 else if (in >= 7961 && in <= 7969) out = 3582;
	 	 	 else if (in >= 7970 && in <= 7978) out = 3583;
	 	 	 else if (in >= 7979 && in <= 7987) out = 3584;
	 	 	 else if (in >= 7988 && in <= 7996) out = 3585;
	 	 	 else if (in >= 7997 && in <= 8006) out = 3586;
	 	 	 else if (in >= 8007 && in <= 8015) out = 3587;
	 	 	 else if (in >= 8016 && in <= 8024) out = 3588;
	 	 	 else if (in >= 8025 && in <= 8033) out = 3589;
	 	 	 else if (in >= 8034 && in <= 8042) out = 3590;
	 	 	 else if (in >= 8043 && in <= 8052) out = 3591;
	 	 	 else if (in >= 8053 && in <= 8061) out = 3592;
	 	 	 else if (in >= 8062 && in <= 8070) out = 3593;
	 	 	 else if (in >= 8071 && in <= 8080) out = 3594;
	 	 	 else if (in >= 8081 && in <= 8089) out = 3595;
	 	 	 else if (in >= 8090 && in <= 8098) out = 3596;
	 	 	 else if (in >= 8099 && in <= 8108) out = 3597;
	 	 	 else if (in >= 8109 && in <= 8117) out = 3598;
	 	 	 else if (in >= 8118 && in <= 8127) out = 3599;
	 	 	 else if (in >= 8128 && in <= 8136) out = 3600;
	 	 	 else if (in >= 8137 && in <= 8145) out = 3601;
	 	 	 else if (in >= 8146 && in <= 8155) out = 3602;
	 	 	 else if (in >= 8156 && in <= 8164) out = 3603;
	 	 	 else if (in >= 8165 && in <= 8174) out = 3604;
	 	 	 else if (in >= 8175 && in <= 8183) out = 3605;
	 	 	 else if (in >= 8184 && in <= 8193) out = 3606;
	 	 	 else if (in >= 8194 && in <= 8202) out = 3607;
	 	 	 else if (in >= 8203 && in <= 8212) out = 3608;
	 	 	 else if (in >= 8213 && in <= 8221) out = 3609;
	 	 	 else if (in >= 8222 && in <= 8231) out = 3610;
	 	 	 else if (in >= 8232 && in <= 8241) out = 3611;
	 	 	 else if (in >= 8242 && in <= 8250) out = 3612;
	 	 	 else if (in >= 8251 && in <= 8260) out = 3613;
	 	 	 else if (in >= 8261 && in <= 8270) out = 3614;
	 	 	 else if (in >= 8271 && in <= 8279) out = 3615;
	 	 	 else if (in >= 8280 && in <= 8289) out = 3616;
	 	 	 else if (in >= 8290 && in <= 8299) out = 3617;
	 	 	 else if (in >= 8300 && in <= 8308) out = 3618;
	 	 	 else if (in >= 8309 && in <= 8318) out = 3619;
	 	 	 else if (in >= 8319 && in <= 8328) out = 3620;
	 	 	 else if (in >= 8329 && in <= 8338) out = 3621;
	 	 	 else if (in >= 8339 && in <= 8347) out = 3622;
	 	 	 else if (in >= 8348 && in <= 8357) out = 3623;
	 	 	 else if (in >= 8358 && in <= 8367) out = 3624;
	 	 	 else if (in >= 8368 && in <= 8377) out = 3625;
	 	 	 else if (in >= 8378 && in <= 8387) out = 3626;
	 	 	 else if (in >= 8388 && in <= 8397) out = 3627;
	 	 	 else if (in >= 8398 && in <= 8407) out = 3628;
	 	 	 else if (in >= 8408 && in <= 8417) out = 3629;
	 	 	 else if (in >= 8418 && in <= 8427) out = 3630;
	 	 	 else if (in >= 8428 && in <= 8436) out = 3631;
	 	 	 else if (in >= 8437 && in <= 8446) out = 3632;
	 	 	 else if (in >= 8447 && in <= 8456) out = 3633;
	 	 	 else if (in >= 8457 && in <= 8466) out = 3634;
	 	 	 else if (in >= 8467 && in <= 8477) out = 3635;
	 	 	 else if (in >= 8478 && in <= 8487) out = 3636;
	 	 	 else if (in >= 8488 && in <= 8497) out = 3637;
	 	 	 else if (in >= 8498 && in <= 8507) out = 3638;
	 	 	 else if (in >= 8508 && in <= 8517) out = 3639;
	 	 	 else if (in >= 8518 && in <= 8527) out = 3640;
	 	 	 else if (in >= 8528 && in <= 8537) out = 3641;
	 	 	 else if (in >= 8538 && in <= 8547) out = 3642;
	 	 	 else if (in >= 8548 && in <= 8558) out = 3643;
	 	 	 else if (in >= 8559 && in <= 8568) out = 3644;
	 	 	 else if (in >= 8569 && in <= 8578) out = 3645;
	 	 	 else if (in >= 8579 && in <= 8588) out = 3646;
	 	 	 else if (in >= 8589 && in <= 8599) out = 3647;
	 	 	 else if (in >= 8600 && in <= 8609) out = 3648;
	 	 	 else if (in >= 8610 && in <= 8619) out = 3649;
	 	 	 else if (in >= 8620 && in <= 8629) out = 3650;
	 	 	 else if (in >= 8630 && in <= 8640) out = 3651;
	 	 	 else if (in >= 8641 && in <= 8650) out = 3652;
	 	 	 else if (in >= 8651 && in <= 8661) out = 3653;
	 	 	 else if (in >= 8662 && in <= 8671) out = 3654;
	 	 	 else if (in >= 8672 && in <= 8681) out = 3655;
	 	 	 else if (in >= 8682 && in <= 8692) out = 3656;
	 	 	 else if (in >= 8693 && in <= 8702) out = 3657;
	 	 	 else if (in >= 8703 && in <= 8713) out = 3658;
	 	 	 else if (in >= 8714 && in <= 8723) out = 3659;
	 	 	 else if (in >= 8724 && in <= 8734) out = 3660;
	 	 	 else if (in >= 8735 && in <= 8745) out = 3661;
	 	 	 else if (in >= 8746 && in <= 8755) out = 3662;
	 	 	 else if (in >= 8756 && in <= 8766) out = 3663;
	 	 	 else if (in >= 8767 && in <= 8776) out = 3664;
	 	 	 else if (in >= 8777 && in <= 8787) out = 3665;
	 	 	 else if (in >= 8788 && in <= 8798) out = 3666;
	 	 	 else if (in >= 8799 && in <= 8808) out = 3667;
	 	 	 else if (in >= 8809 && in <= 8819) out = 3668;
	 	 	 else if (in >= 8820 && in <= 8830) out = 3669;
	 	 	 else if (in >= 8831 && in <= 8841) out = 3670;
	 	 	 else if (in >= 8842 && in <= 8851) out = 3671;
	 	 	 else if (in >= 8852 && in <= 8862) out = 3672;
	 	 	 else if (in >= 8863 && in <= 8873) out = 3673;
	 	 	 else if (in >= 8874 && in <= 8884) out = 3674;
	 	 	 else if (in >= 8885 && in <= 8895) out = 3675;
	 	 	 else if (in >= 8896 && in <= 8906) out = 3676;
	 	 	 else if (in >= 8907 && in <= 8917) out = 3677;
	 	 	 else if (in >= 8918 && in <= 8928) out = 3678;
	 	 	 else if (in >= 8929 && in <= 8939) out = 3679;
	 	 	 else if (in >= 8940 && in <= 8950) out = 3680;
	 	 	 else if (in >= 8951 && in <= 8961) out = 3681;
	 	 	 else if (in >= 8962 && in <= 8972) out = 3682;
	 	 	 else if (in >= 8973 && in <= 8983) out = 3683;
	 	 	 else if (in >= 8984 && in <= 8994) out = 3684;
	 	 	 else if (in >= 8995 && in <= 9005) out = 3685;
	 	 	 else if (in >= 9006 && in <= 9016) out = 3686;
	 	 	 else if (in >= 9017 && in <= 9027) out = 3687;
	 	 	 else if (in >= 9028 && in <= 9038) out = 3688;
	 	 	 else if (in >= 9039 && in <= 9050) out = 3689;
	 	 	 else if (in >= 9051 && in <= 9061) out = 3690;
	 	 	 else if (in >= 9062 && in <= 9072) out = 3691;
	 	 	 else if (in >= 9073 && in <= 9083) out = 3692;
	 	 	 else if (in >= 9084 && in <= 9095) out = 3693;
	 	 	 else if (in >= 9096 && in <= 9106) out = 3694;
	 	 	 else if (in >= 9107 && in <= 9117) out = 3695;
	 	 	 else if (in >= 9118 && in <= 9129) out = 3696;
	 	 	 else if (in >= 9130 && in <= 9140) out = 3697;
	 	 	 else if (in >= 9141 && in <= 9152) out = 3698;
	 	 	 else if (in >= 9153 && in <= 9163) out = 3699;
	 	 	 else if (in >= 9164 && in <= 9175) out = 3700;
	 	 	 else if (in >= 9176 && in <= 9186) out = 3701;
	 	 	 else if (in >= 9187 && in <= 9198) out = 3702;
	 	 	 else if (in >= 9199 && in <= 9209) out = 3703;
	 	 	 else if (in >= 9210 && in <= 9221) out = 3704;
	 	 	 else if (in >= 9222 && in <= 9232) out = 3705;
	 	 	 else if (in >= 9233 && in <= 9244) out = 3706;
	 	 	 else if (in >= 9245 && in <= 9256) out = 3707;
	 	 	 else if (in >= 9257 && in <= 9267) out = 3708;
	 	 	 else if (in >= 9268 && in <= 9279) out = 3709;
	 	 	 else if (in >= 9280 && in <= 9291) out = 3710;
	 	 	 else if (in >= 9292 && in <= 9303) out = 3711;
	 	 	 else if (in >= 9304 && in <= 9315) out = 3712;
	 	 	 else if (in >= 9316 && in <= 9326) out = 3713;
	 	 	 else if (in >= 9327 && in <= 9338) out = 3714;
	 	 	 else if (in >= 9339 && in <= 9350) out = 3715;
	 	 	 else if (in >= 9351 && in <= 9362) out = 3716;
	 	 	 else if (in >= 9363 && in <= 9374) out = 3717;
	 	 	 else if (in >= 9375 && in <= 9386) out = 3718;
	 	 	 else if (in >= 9387 && in <= 9398) out = 3719;
	 	 	 else if (in >= 9399 && in <= 9410) out = 3720;
	 	 	 else if (in >= 9411 && in <= 9422) out = 3721;
	 	 	 else if (in >= 9423 && in <= 9434) out = 3722;
	 	 	 else if (in >= 9435 && in <= 9446) out = 3723;
	 	 	 else if (in >= 9447 && in <= 9458) out = 3724;
	 	 	 else if (in >= 9459 && in <= 9471) out = 3725;
	 	 	 else if (in >= 9472 && in <= 9483) out = 3726;
	 	 	 else if (in >= 9484 && in <= 9495) out = 3727;
	 	 	 else if (in >= 9496 && in <= 9507) out = 3728;
	 	 	 else if (in >= 9508 && in <= 9520) out = 3729;
	 	 	 else if (in >= 9521 && in <= 9532) out = 3730;
	 	 	 else if (in >= 9533 && in <= 9544) out = 3731;
	 	 	 else if (in >= 9545 && in <= 9557) out = 3732;
	 	 	 else if (in >= 9558 && in <= 9569) out = 3733;
	 	 	 else if (in >= 9570 && in <= 9582) out = 3734;
	 	 	 else if (in >= 9583 && in <= 9594) out = 3735;
	 	 	 else if (in >= 9595 && in <= 9607) out = 3736;
	 	 	 else if (in >= 9608 && in <= 9619) out = 3737;
	 	 	 else if (in >= 9620 && in <= 9632) out = 3738;
	 	 	 else if (in >= 9633 && in <= 9644) out = 3739;
	 	 	 else if (in >= 9645 && in <= 9657) out = 3740;
	 	 	 else if (in >= 9658 && in <= 9670) out = 3741;
	 	 	 else if (in >= 9671 && in <= 9682) out = 3742;
	 	 	 else if (in >= 9683 && in <= 9695) out = 3743;
	 	 	 else if (in >= 9696 && in <= 9708) out = 3744;
	 	 	 else if (in >= 9709 && in <= 9721) out = 3745;
	 	 	 else if (in >= 9722 && in <= 9734) out = 3746;
	 	 	 else if (in >= 9735 && in <= 9747) out = 3747;
	 	 	 else if (in >= 9748 && in <= 9759) out = 3748;
	 	 	 else if (in >= 9760 && in <= 9772) out = 3749;
	 	 	 else if (in >= 9773 && in <= 9785) out = 3750;
	 	 	 else if (in >= 9786 && in <= 9798) out = 3751;
	 	 	 else if (in >= 9799 && in <= 9811) out = 3752;
	 	 	 else if (in >= 9812 && in <= 9825) out = 3753;
	 	 	 else if (in >= 9826 && in <= 9838) out = 3754;
	 	 	 else if (in >= 9839 && in <= 9851) out = 3755;
	 	 	 else if (in >= 9852 && in <= 9864) out = 3756;
	 	 	 else if (in >= 9865 && in <= 9877) out = 3757;
	 	 	 else if (in >= 9878 && in <= 9891) out = 3758;
	 	 	 else if (in >= 9892 && in <= 9904) out = 3759;
	 	 	 else if (in >= 9905 && in <= 9917) out = 3760;
	 	 	 else if (in >= 9918 && in <= 9931) out = 3761;
	 	 	 else if (in >= 9932 && in <= 9944) out = 3762;
	 	 	 else if (in >= 9945 && in <= 9957) out = 3763;
	 	 	 else if (in >= 9958 && in <= 9971) out = 3764;
	 	 	 else if (in >= 9972 && in <= 9984) out = 3765;
	 	 	 else if (in >= 9985 && in <= 9998) out = 3766;
	 	 	 else if (in >= 9999 && in <= 10012) out = 3767;
	 	 	 else if (in >= 10013 && in <= 10025) out = 3768;
	 	 	 else if (in >= 10026 && in <= 10039) out = 3769;
	 	 	 else if (in >= 10040 && in <= 10053) out = 3770;
	 	 	 else if (in >= 10054 && in <= 10066) out = 3771;
	 	 	 else if (in >= 10067 && in <= 10080) out = 3772;
	 	 	 else if (in >= 10081 && in <= 10094) out = 3773;
	 	 	 else if (in >= 10095 && in <= 10108) out = 3774;
	 	 	 else if (in >= 10109 && in <= 10122) out = 3775;
	 	 	 else if (in >= 10123 && in <= 10136) out = 3776;
	 	 	 else if (in >= 10137 && in <= 10150) out = 3777;
	 	 	 else if (in >= 10151 && in <= 10164) out = 3778;
	 	 	 else if (in >= 10165 && in <= 10178) out = 3779;
	 	 	 else if (in >= 10179 && in <= 10192) out = 3780;
	 	 	 else if (in >= 10193 && in <= 10206) out = 3781;
	 	 	 else if (in >= 10207 && in <= 10220) out = 3782;
	 	 	 else if (in >= 10221 && in <= 10234) out = 3783;
	 	 	 else if (in >= 10235 && in <= 10249) out = 3784;
	 	 	 else if (in >= 10250 && in <= 10263) out = 3785;
	 	 	 else if (in >= 10264 && in <= 10277) out = 3786;
	 	 	 else if (in >= 10278 && in <= 10292) out = 3787;
	 	 	 else if (in >= 10293 && in <= 10306) out = 3788;
	 	 	 else if (in >= 10307 && in <= 10321) out = 3789;
	 	 	 else if (in >= 10322 && in <= 10335) out = 3790;
	 	 	 else if (in >= 10336 && in <= 10350) out = 3791;
	 	 	 else if (in >= 10351 && in <= 10364) out = 3792;
	 	 	 else if (in >= 10365 && in <= 10379) out = 3793;
	 	 	 else if (in >= 10380 && in <= 10394) out = 3794;
	 	 	 else if (in >= 10395 && in <= 10408) out = 3795;
	 	 	 else if (in >= 10409 && in <= 10423) out = 3796;
	 	 	 else if (in >= 10424 && in <= 10438) out = 3797;
	 	 	 else if (in >= 10439 && in <= 10453) out = 3798;
	 	 	 else if (in >= 10454 && in <= 10468) out = 3799;
	 	 	 else if (in >= 10469 && in <= 10483) out = 3800;
	 	 	 else if (in >= 10484 && in <= 10498) out = 3801;
	 	 	 else if (in >= 10499 && in <= 10513) out = 3802;
	 	 	 else if (in >= 10514 && in <= 10528) out = 3803;
	 	 	 else if (in >= 10529 && in <= 10543) out = 3804;
	 	 	 else if (in >= 10544 && in <= 10559) out = 3805;
	 	 	 else if (in >= 10560 && in <= 10574) out = 3806;
	 	 	 else if (in >= 10575 && in <= 10589) out = 3807;
	 	 	 else if (in >= 10590 && in <= 10605) out = 3808;
	 	 	 else if (in >= 10606 && in <= 10620) out = 3809;
	 	 	 else if (in >= 10621 && in <= 10635) out = 3810;
	 	 	 else if (in >= 10636 && in <= 10651) out = 3811;
	 	 	 else if (in >= 10652 && in <= 10667) out = 3812;
	 	 	 else if (in >= 10668 && in <= 10682) out = 3813;
	 	 	 else if (in >= 10683 && in <= 10698) out = 3814;
	 	 	 else if (in >= 10699 && in <= 10714) out = 3815;
	 	 	 else if (in >= 10715 && in <= 10729) out = 3816;
	 	 	 else if (in >= 10730 && in <= 10745) out = 3817;
	 	 	 else if (in >= 10746 && in <= 10761) out = 3818;
	 	 	 else if (in >= 10762 && in <= 10777) out = 3819;
	 	 	 else if (in >= 10778 && in <= 10793) out = 3820;
	 	 	 else if (in >= 10794 && in <= 10809) out = 3821;
	 	 	 else if (in >= 10810 && in <= 10825) out = 3822;
	 	 	 else if (in >= 10826 && in <= 10841) out = 3823;
	 	 	 else if (in >= 10842 && in <= 10858) out = 3824;
	 	 	 else if (in >= 10859 && in <= 10874) out = 3825;
	 	 	 else if (in >= 10875 && in <= 10890) out = 3826;
	 	 	 else if (in >= 10891 && in <= 10907) out = 3827;
	 	 	 else if (in >= 10908 && in <= 10923) out = 3828;
	 	 	 else if (in >= 10924 && in <= 10939) out = 3829;
	 	 	 else if (in >= 10940 && in <= 10956) out = 3830;
	 	 	 else if (in >= 10957 && in <= 10973) out = 3831;
	 	 	 else if (in >= 10974 && in <= 10989) out = 3832;
	 	 	 else if (in >= 10990 && in <= 11006) out = 3833;
	 	 	 else if (in >= 11007 && in <= 11023) out = 3834;
	 	 	 else if (in >= 11024 && in <= 11040) out = 3835;
	 	 	 else if (in >= 11041 && in <= 11057) out = 3836;
	 	 	 else if (in >= 11058 && in <= 11074) out = 3837;
	 	 	 else if (in >= 11075 && in <= 11091) out = 3838;
	 	 	 else if (in >= 11092 && in <= 11108) out = 3839;
	 	 	 else if (in >= 11109 && in <= 11125) out = 3840;
	 	 	 else if (in >= 11126 && in <= 11142) out = 3841;
	 	 	 else if (in >= 11143 && in <= 11159) out = 3842;
	 	 	 else if (in >= 11160 && in <= 11177) out = 3843;
	 	 	 else if (in >= 11178 && in <= 11194) out = 3844;
	 	 	 else if (in >= 11195 && in <= 11212) out = 3845;
	 	 	 else if (in >= 11213 && in <= 11229) out = 3846;
	 	 	 else if (in >= 11230 && in <= 11247) out = 3847;
	 	 	 else if (in >= 11248 && in <= 11264) out = 3848;
	 	 	 else if (in >= 11265 && in <= 11282) out = 3849;
	 	 	 else if (in >= 11283 && in <= 11300) out = 3850;
	 	 	 else if (in >= 11301 && in <= 11318) out = 3851;
	 	 	 else if (in >= 11319 && in <= 11336) out = 3852;
	 	 	 else if (in >= 11337 && in <= 11354) out = 3853;
	 	 	 else if (in >= 11355 && in <= 11372) out = 3854;
	 	 	 else if (in >= 11373 && in <= 11390) out = 3855;
	 	 	 else if (in >= 11391 && in <= 11408) out = 3856;
	 	 	 else if (in >= 11409 && in <= 11427) out = 3857;
	 	 	 else if (in >= 11428 && in <= 11445) out = 3858;
	 	 	 else if (in >= 11446 && in <= 11464) out = 3859;
	 	 	 else if (in >= 11465 && in <= 11482) out = 3860;
	 	 	 else if (in >= 11483 && in <= 11501) out = 3861;
	 	 	 else if (in >= 11502 && in <= 11519) out = 3862;
	 	 	 else if (in >= 11520 && in <= 11538) out = 3863;
	 	 	 else if (in >= 11539 && in <= 11557) out = 3864;
	 	 	 else if (in >= 11558 && in <= 11576) out = 3865;
	 	 	 else if (in >= 11577 && in <= 11595) out = 3866;
	 	 	 else if (in >= 11596 && in <= 11614) out = 3867;
	 	 	 else if (in >= 11615 && in <= 11633) out = 3868;
	 	 	 else if (in >= 11634 && in <= 11652) out = 3869;
	 	 	 else if (in >= 11653 && in <= 11672) out = 3870;
	 	 	 else if (in >= 11673 && in <= 11691) out = 3871;
	 	 	 else if (in >= 11692 && in <= 11710) out = 3872;
	 	 	 else if (in >= 11711 && in <= 11730) out = 3873;
	 	 	 else if (in >= 11731 && in <= 11750) out = 3874;
	 	 	 else if (in >= 11751 && in <= 11769) out = 3875;
	 	 	 else if (in >= 11770 && in <= 11789) out = 3876;
	 	 	 else if (in >= 11790 && in <= 11809) out = 3877;
	 	 	 else if (in >= 11810 && in <= 11829) out = 3878;
	 	 	 else if (in >= 11830 && in <= 11849) out = 3879;
	 	 	 else if (in >= 11850 && in <= 11869) out = 3880;
	 	 	 else if (in >= 11870 && in <= 11889) out = 3881;
	 	 	 else if (in >= 11890 && in <= 11910) out = 3882;
	 	 	 else if (in >= 11911 && in <= 11930) out = 3883;
	 	 	 else if (in >= 11931 && in <= 11951) out = 3884;
	 	 	 else if (in >= 11952 && in <= 11971) out = 3885;
	 	 	 else if (in >= 11972 && in <= 11992) out = 3886;
	 	 	 else if (in >= 11993 && in <= 12013) out = 3887;
	 	 	 else if (in >= 12014 && in <= 12034) out = 3888;
	 	 	 else if (in >= 12035 && in <= 12055) out = 3889;
	 	 	 else if (in >= 12056 && in <= 12076) out = 3890;
	 	 	 else if (in >= 12077 && in <= 12097) out = 3891;
	 	 	 else if (in >= 12098 && in <= 12118) out = 3892;
	 	 	 else if (in >= 12119 && in <= 12140) out = 3893;
	 	 	 else if (in >= 12141 && in <= 12161) out = 3894;
	 	 	 else if (in >= 12162 && in <= 12183) out = 3895;
	 	 	 else if (in >= 12184 && in <= 12204) out = 3896;
	 	 	 else if (in >= 12205 && in <= 12226) out = 3897;
	 	 	 else if (in >= 12227 && in <= 12248) out = 3898;
	 	 	 else if (in >= 12249 && in <= 12270) out = 3899;
	 	 	 else if (in >= 12271 && in <= 12292) out = 3900;
	 	 	 else if (in >= 12293 && in <= 12314) out = 3901;
	 	 	 else if (in >= 12315 && in <= 12337) out = 3902;
	 	 	 else if (in >= 12338 && in <= 12359) out = 3903;
	 	 	 else if (in >= 12360 && in <= 12382) out = 3904;
	 	 	 else if (in >= 12383 && in <= 12404) out = 3905;
	 	 	 else if (in >= 12405 && in <= 12427) out = 3906;
	 	 	 else if (in >= 12428 && in <= 12450) out = 3907;
	 	 	 else if (in >= 12451 && in <= 12473) out = 3908;
	 	 	 else if (in >= 12474 && in <= 12496) out = 3909;
	 	 	 else if (in >= 12497 && in <= 12519) out = 3910;
	 	 	 else if (in >= 12520 && in <= 12543) out = 3911;
	 	 	 else if (in >= 12544 && in <= 12566) out = 3912;
	 	 	 else if (in >= 12567 && in <= 12590) out = 3913;
	 	 	 else if (in >= 12591 && in <= 12614) out = 3914;
	 	 	 else if (in >= 12615 && in <= 12637) out = 3915;
	 	 	 else if (in >= 12638 && in <= 12661) out = 3916;
	 	 	 else if (in >= 12662 && in <= 12686) out = 3917;
	 	 	 else if (in >= 12687 && in <= 12710) out = 3918;
	 	 	 else if (in >= 12711 && in <= 12734) out = 3919;
	 	 	 else if (in >= 12735 && in <= 12759) out = 3920;
	 	 	 else if (in >= 12760 && in <= 12783) out = 3921;
	 	 	 else if (in >= 12784 && in <= 12808) out = 3922;
	 	 	 else if (in >= 12809 && in <= 12833) out = 3923;
	 	 	 else if (in >= 12834 && in <= 12858) out = 3924;
	 	 	 else if (in >= 12859 && in <= 12883) out = 3925;
	 	 	 else if (in >= 12884 && in <= 12909) out = 3926;
	 	 	 else if (in >= 12910 && in <= 12934) out = 3927;
	 	 	 else if (in >= 12935 && in <= 12960) out = 3928;
	 	 	 else if (in >= 12961 && in <= 12986) out = 3929;
	 	 	 else if (in >= 12987 && in <= 13012) out = 3930;
	 	 	 else if (in >= 13013 && in <= 13038) out = 3931;
	 	 	 else if (in >= 13039 && in <= 13064) out = 3932;
	 	 	 else if (in >= 13065 && in <= 13090) out = 3933;
	 	 	 else if (in >= 13091 && in <= 13117) out = 3934;
	 	 	 else if (in >= 13118 && in <= 13144) out = 3935;
	 	 	 else if (in >= 13145 && in <= 13171) out = 3936;
	 	 	 else if (in >= 13172 && in <= 13198) out = 3937;
	 	 	 else if (in >= 13199 && in <= 13225) out = 3938;
	 	 	 else if (in >= 13226 && in <= 13252) out = 3939;
	 	 	 else if (in >= 13253 && in <= 13280) out = 3940;
	 	 	 else if (in >= 13281 && in <= 13307) out = 3941;
	 	 	 else if (in >= 13308 && in <= 13335) out = 3942;
	 	 	 else if (in >= 13336 && in <= 13363) out = 3943;
	 	 	 else if (in >= 13364 && in <= 13392) out = 3944;
	 	 	 else if (in >= 13393 && in <= 13420) out = 3945;
	 	 	 else if (in >= 13421 && in <= 13449) out = 3946;
	 	 	 else if (in >= 13450 && in <= 13478) out = 3947;
	 	 	 else if (in >= 13479 && in <= 13507) out = 3948;
	 	 	 else if (in >= 13508 && in <= 13536) out = 3949;
	 	 	 else if (in >= 13537 && in <= 13565) out = 3950;
	 	 	 else if (in >= 13566 && in <= 13595) out = 3951;
	 	 	 else if (in >= 13596 && in <= 13624) out = 3952;
	 	 	 else if (in >= 13625 && in <= 13654) out = 3953;
	 	 	 else if (in >= 13655 && in <= 13685) out = 3954;
	 	 	 else if (in >= 13686 && in <= 13715) out = 3955;
	 	 	 else if (in >= 13716 && in <= 13746) out = 3956;
	 	 	 else if (in >= 13747 && in <= 13776) out = 3957;
	 	 	 else if (in >= 13777 && in <= 13807) out = 3958;
	 	 	 else if (in >= 13808 && in <= 13839) out = 3959;
	 	 	 else if (in >= 13840 && in <= 13870) out = 3960;
	 	 	 else if (in >= 13871 && in <= 13902) out = 3961;
	 	 	 else if (in >= 13903 && in <= 13934) out = 3962;
	 	 	 else if (in >= 13935 && in <= 13966) out = 3963;
	 	 	 else if (in >= 13967 && in <= 13999) out = 3964;
	 	 	 else if (in >= 14000 && in <= 14031) out = 3965;
	 	 	 else if (in >= 14032 && in <= 14064) out = 3966;
	 	 	 else if (in >= 14065 && in <= 14097) out = 3967;
	 	 	 else if (in >= 14098 && in <= 14131) out = 3968;
	 	 	 else if (in >= 14132 && in <= 14164) out = 3969;
	 	 	 else if (in >= 14165 && in <= 14198) out = 3970;
	 	 	 else if (in >= 14199 && in <= 14232) out = 3971;
	 	 	 else if (in >= 14233 && in <= 14267) out = 3972;
	 	 	 else if (in >= 14268 && in <= 14302) out = 3973;
	 	 	 else if (in >= 14303 && in <= 14337) out = 3974;
	 	 	 else if (in >= 14338 && in <= 14372) out = 3975;
	 	 	 else if (in >= 14373 && in <= 14408) out = 3976;
	 	 	 else if (in >= 14409 && in <= 14443) out = 3977;
	 	 	 else if (in >= 14444 && in <= 14480) out = 3978;
	 	 	 else if (in >= 14481 && in <= 14516) out = 3979;
	 	 	 else if (in >= 14517 && in <= 14553) out = 3980;
	 	 	 else if (in >= 14554 && in <= 14590) out = 3981;
	 	 	 else if (in >= 14591 && in <= 14628) out = 3982;
	 	 	 else if (in >= 14629 && in <= 14665) out = 3983;
	 	 	 else if (in >= 14666 && in <= 14703) out = 3984;
	 	 	 else if (in >= 14704 && in <= 14742) out = 3985;
	 	 	 else if (in >= 14743 && in <= 14781) out = 3986;
	 	 	 else if (in >= 14782 && in <= 14820) out = 3987;
	 	 	 else if (in >= 14821 && in <= 14859) out = 3988;
	 	 	 else if (in >= 14860 && in <= 14899) out = 3989;
	 	 	 else if (in >= 14900 && in <= 14939) out = 3990;
	 	 	 else if (in >= 14940 && in <= 14980) out = 3991;
	 	 	 else if (in >= 14981 && in <= 15021) out = 3992;
	 	 	 else if (in >= 15022 && in <= 15062) out = 3993;
	 	 	 else if (in >= 15063 && in <= 15104) out = 3994;
	 	 	 else if (in >= 15105 && in <= 15146) out = 3995;
	 	 	 else if (in >= 15147 && in <= 15189) out = 3996;
	 	 	 else if (in >= 15190 && in <= 15232) out = 3997;
	 	 	 else if (in >= 15233 && in <= 15275) out = 3998;
	 	 	 else if (in >= 15276 && in <= 15319) out = 3999;
	 	 	 else if (in >= 15320 && in <= 15364) out = 4000;
	 	 	 else if (in >= 15365 && in <= 15408) out = 4001;
	 	 	 else if (in >= 15409 && in <= 15454) out = 4002;
	 	 	 else if (in >= 15455 && in <= 15500) out = 4003;
	 	 	 else if (in >= 15501 && in <= 15546) out = 4004;
	 	 	 else if (in >= 15547 && in <= 15593) out = 4005;
	 	 	 else if (in >= 15594 && in <= 15640) out = 4006;
	 	 	 else if (in >= 15641 && in <= 15688) out = 4007;
	 	 	 else if (in >= 15689 && in <= 15736) out = 4008;
	 	 	 else if (in >= 15737 && in <= 15785) out = 4009;
	 	 	 else if (in >= 15786 && in <= 15835) out = 4010;
	 	 	 else if (in >= 15836 && in <= 15885) out = 4011;
	 	 	 else if (in >= 15886 && in <= 15935) out = 4012;
	 	 	 else if (in >= 15936 && in <= 15987) out = 4013;
	 	 	 else if (in >= 15988 && in <= 16038) out = 4014;
	 	 	 else if (in >= 16039 && in <= 16091) out = 4015;
	 	 	 else if (in >= 16092 && in <= 16144) out = 4016;
	 	 	 else if (in >= 16145 && in <= 16198) out = 4017;
	 	 	 else if (in >= 16199 && in <= 16253) out = 4018;
	 	 	 else if (in >= 16254 && in <= 16308) out = 4019;
	 	 	 else if (in >= 16309 && in <= 16364) out = 4020;
	 	 	 else if (in >= 16365 && in <= 16421) out = 4021;
	 	 	 else if (in >= 16422 && in <= 16478) out = 4022;
	 	 	 else if (in >= 16479 && in <= 16536) out = 4023;
	 	 	 else if (in >= 16537 && in <= 16596) out = 4024;
	 	 	 else if (in >= 16597 && in <= 16656) out = 4025;
	 	 	 else if (in >= 16657 && in <= 16716) out = 4026;
	 	 	 else if (in >= 16717 && in <= 16778) out = 4027;
	 	 	 else if (in >= 16779 && in <= 16841) out = 4028;
	 	 	 else if (in >= 16842 && in <= 16904) out = 4029;
	 	 	 else if (in >= 16905 && in <= 16969) out = 4030;
	 	 	 else if (in >= 16970 && in <= 17034) out = 4031;
	 	 	 else if (in >= 17035 && in <= 17101) out = 4032;
	 	 	 else if (in >= 17102 && in <= 17168) out = 4033;
	 	 	 else if (in >= 17169 && in <= 17237) out = 4034;
	 	 	 else if (in >= 17238 && in <= 17307) out = 4035;
	 	 	 else if (in >= 17308 && in <= 17378) out = 4036;
	 	 	 else if (in >= 17379 && in <= 17450) out = 4037;
	 	 	 else if (in >= 17451 && in <= 17524) out = 4038;
	 	 	 else if (in >= 17525 && in <= 17599) out = 4039;
	 	 	 else if (in >= 17600 && in <= 17675) out = 4040;
	 	 	 else if (in >= 17676 && in <= 17752) out = 4041;
	 	 	 else if (in >= 17753 && in <= 17831) out = 4042;
	 	 	 else if (in >= 17832 && in <= 17912) out = 4043;
	 	 	 else if (in >= 17913 && in <= 17994) out = 4044;
	 	 	 else if (in >= 17995 && in <= 18078) out = 4045;
	 	 	 else if (in >= 18079 && in <= 18163) out = 4046;
	 	 	 else if (in >= 18164 && in <= 18251) out = 4047;
	 	 	 else if (in >= 18252 && in <= 18340) out = 4048;
	 	 	 else if (in >= 18341 && in <= 18431) out = 4049;
	 	 	 else if (in >= 18432 && in <= 18524) out = 4050;
	 	 	 else if (in >= 18525 && in <= 18619) out = 4051;
	 	 	 else if (in >= 18620 && in <= 18716) out = 4052;
	 	 	 else if (in >= 18717 && in <= 18816) out = 4053;
	 	 	 else if (in >= 18817 && in <= 18918) out = 4054;
	 	 	 else if (in >= 18919 && in <= 19023) out = 4055;
	 	 	 else if (in >= 19024 && in <= 19130) out = 4056;
	 	 	 else if (in >= 19131 && in <= 19241) out = 4057;
	 	 	 else if (in >= 19242 && in <= 19354) out = 4058;
	 	 	 else if (in >= 19355 && in <= 19470) out = 4059;
	 	 	 else if (in >= 19471 && in <= 19590) out = 4060;
	 	 	 else if (in >= 19591 && in <= 19713) out = 4061;
	 	 	 else if (in >= 19714 && in <= 19840) out = 4062;
	 	 	 else if (in >= 19841 && in <= 19971) out = 4063;
	 	 	 else if (in >= 19972 && in <= 20107) out = 4064;
	 	 	 else if (in >= 20108 && in <= 20247) out = 4065;
	 	 	 else if (in >= 20248 && in <= 20391) out = 4066;
	 	 	 else if (in >= 20392 && in <= 20541) out = 4067;
	 	 	 else if (in >= 20542 && in <= 20697) out = 4068;
	 	 	 else if (in >= 20698 && in <= 20858) out = 4069;
	 	 	 else if (in >= 20859 && in <= 21027) out = 4070;
	 	 	 else if (in >= 21028 && in <= 21202) out = 4071;
	 	 	 else if (in >= 21203 && in <= 21385) out = 4072;
	 	 	 else if (in >= 21386 && in <= 21577) out = 4073;
	 	 	 else if (in >= 21578 && in <= 21777) out = 4074;
	 	 	 else if (in >= 21778 && in <= 21989) out = 4075;
	 	 	 else if (in >= 21990 && in <= 22211) out = 4076;
	 	 	 else if (in >= 22212 && in <= 22446) out = 4077;
	 	 	 else if (in >= 22447 && in <= 22696) out = 4078;
	 	 	 else if (in >= 22697 && in <= 22961) out = 4079;
	 	 	 else if (in >= 22962 && in <= 23244) out = 4080;
	 	 	 else if (in >= 23245 && in <= 23549) out = 4081;
	 	 	 else if (in >= 23550 && in <= 23878) out = 4082;
	 	 	 else if (in >= 23879 && in <= 24235) out = 4083;
	 	 	 else if (in >= 24236 && in <= 24627) out = 4084;
	 	 	 else if (in >= 24628 && in <= 25059) out = 4085;
	 	 	 else if (in >= 25060 && in <= 25543) out = 4086;
	 	 	 else if (in >= 25544 && in <= 26091) out = 4087;
	 	 	 else if (in >= 26092 && in <= 26723) out = 4088;
	 	 	 else if (in >= 26724 && in <= 27471) out = 4089;
	 	 	 else if (in >= 27472 && in <= 28386) out = 4090;
	 	 	 else if (in >= 28387 && in <= 29565) out = 4091;
	 	 	 else if (in >= 29566 && in <= 31227) out = 4092;
	 	 	 else if (in >= 31228 && in <= 34067) out = 4093;
	 	 	 else if (in >= 34068 && in <= 65535) out = 4094;
	 	 	else out=4095;
	 endmodule
	 
	 
module log_int(input logic [12:0] in,
	 output logic [16:0] out);
	 	 always_comb
	 	 	 if (in == 0) out = -66019;
	 	 	 else if (in == 1) out = -34069;
	 	 	 else if (in == 2) out = -31230;
	 	 	 else if (in == 3) out = -29569;
	 	 	 else if (in == 4) out = -28391;
	 	 	 else if (in == 5) out = -27477;
	 	 	 else if (in == 6) out = -26730;
	 	 	 else if (in == 7) out = -26099;
	 	 	 else if (in == 8) out = -25552;
	 	 	 else if (in == 9) out = -25069;
	 	 	 else if (in == 10) out = -24638;
	 	 	 else if (in == 11) out = -24247;
	 	 	 else if (in == 12) out = -23891;
	 	 	 else if (in == 13) out = -23563;
	 	 	 else if (in == 14) out = -23259;
	 	 	 else if (in == 15) out = -22977;
	 	 	 else if (in == 16) out = -22713;
	 	 	 else if (in == 17) out = -22464;
	 	 	 else if (in == 18) out = -22230;
	 	 	 else if (in == 19) out = -22009;
	 	 	 else if (in == 20) out = -21799;
	 	 	 else if (in == 21) out = -21599;
	 	 	 else if (in == 22) out = -21408;
	 	 	 else if (in == 23) out = -21226;
	 	 	 else if (in == 24) out = -21052;
	 	 	 else if (in == 25) out = -20885;
	 	 	 else if (in == 26) out = -20724;
	 	 	 else if (in == 27) out = -20569;
	 	 	 else if (in == 28) out = -20420;
	 	 	 else if (in == 29) out = -20277;
	 	 	 else if (in == 30) out = -20138;
	 	 	 else if (in == 31) out = -20003;
	 	 	 else if (in == 32) out = -19873;
	 	 	 else if (in == 33) out = -19747;
	 	 	 else if (in == 34) out = -19625;
	 	 	 else if (in == 35) out = -19506;
	 	 	 else if (in == 36) out = -19391;
	 	 	 else if (in == 37) out = -19279;
	 	 	 else if (in == 38) out = -19170;
	 	 	 else if (in == 39) out = -19063;
	 	 	 else if (in == 40) out = -18959;
	 	 	 else if (in == 41) out = -18858;
	 	 	 else if (in == 42) out = -18760;
	 	 	 else if (in == 43) out = -18663;
	 	 	 else if (in == 44) out = -18569;
	 	 	 else if (in == 45) out = -18477;
	 	 	 else if (in == 46) out = -18387;
	 	 	 else if (in == 47) out = -18299;
	 	 	 else if (in == 48) out = -18213;
	 	 	 else if (in == 49) out = -18128;
	 	 	 else if (in == 50) out = -18045;
	 	 	 else if (in == 51) out = -17964;
	 	 	 else if (in == 52) out = -17885;
	 	 	 else if (in == 53) out = -17807;
	 	 	 else if (in == 54) out = -17730;
	 	 	 else if (in == 55) out = -17655;
	 	 	 else if (in == 56) out = -17581;
	 	 	 else if (in == 57) out = -17509;
	 	 	 else if (in == 58) out = -17437;
	 	 	 else if (in == 59) out = -17367;
	 	 	 else if (in == 60) out = -17299;
	 	 	 else if (in == 61) out = -17231;
	 	 	 else if (in == 62) out = -17164;
	 	 	 else if (in == 63) out = -17099;
	 	 	 else if (in == 64) out = -17034;
	 	 	 else if (in == 65) out = -16971;
	 	 	 else if (in == 66) out = -16908;
	 	 	 else if (in == 67) out = -16847;
	 	 	 else if (in == 68) out = -16786;
	 	 	 else if (in == 69) out = -16726;
	 	 	 else if (in == 70) out = -16667;
	 	 	 else if (in == 71) out = -16609;
	 	 	 else if (in == 72) out = -16552;
	 	 	 else if (in == 73) out = -16495;
	 	 	 else if (in == 74) out = -16440;
	 	 	 else if (in == 75) out = -16385;
	 	 	 else if (in == 76) out = -16330;
	 	 	 else if (in == 77) out = -16277;
	 	 	 else if (in == 78) out = -16224;
	 	 	 else if (in == 79) out = -16172;
	 	 	 else if (in == 80) out = -16120;
	 	 	 else if (in == 81) out = -16069;
	 	 	 else if (in == 82) out = -16019;
	 	 	 else if (in == 83) out = -15969;
	 	 	 else if (in == 84) out = -15920;
	 	 	 else if (in == 85) out = -15872;
	 	 	 else if (in == 86) out = -15824;
	 	 	 else if (in == 87) out = -15777;
	 	 	 else if (in == 88) out = -15730;
	 	 	 else if (in == 89) out = -15684;
	 	 	 else if (in == 90) out = -15638;
	 	 	 else if (in == 91) out = -15593;
	 	 	 else if (in == 92) out = -15548;
	 	 	 else if (in == 93) out = -15504;
	 	 	 else if (in == 94) out = -15460;
	 	 	 else if (in == 95) out = -15416;
	 	 	 else if (in == 96) out = -15374;
	 	 	 else if (in == 97) out = -15331;
	 	 	 else if (in == 98) out = -15289;
	 	 	 else if (in == 99) out = -15247;
	 	 	 else if (in == 100) out = -15206;
	 	 	 else if (in == 101) out = -15166;
	 	 	 else if (in == 102) out = -15125;
	 	 	 else if (in == 103) out = -15085;
	 	 	 else if (in == 104) out = -15046;
	 	 	 else if (in == 105) out = -15006;
	 	 	 else if (in == 106) out = -14968;
	 	 	 else if (in == 107) out = -14929;
	 	 	 else if (in == 108) out = -14891;
	 	 	 else if (in == 109) out = -14853;
	 	 	 else if (in == 110) out = -14816;
	 	 	 else if (in == 111) out = -14779;
	 	 	 else if (in == 112) out = -14742;
	 	 	 else if (in == 113) out = -14706;
	 	 	 else if (in == 114) out = -14670;
	 	 	 else if (in == 115) out = -14634;
	 	 	 else if (in == 116) out = -14598;
	 	 	 else if (in == 117) out = -14563;
	 	 	 else if (in == 118) out = -14528;
	 	 	 else if (in == 119) out = -14494;
	 	 	 else if (in == 120) out = -14460;
	 	 	 else if (in == 121) out = -14426;
	 	 	 else if (in == 122) out = -14392;
	 	 	 else if (in == 123) out = -14358;
	 	 	 else if (in == 124) out = -14325;
	 	 	 else if (in == 125) out = -14292;
	 	 	 else if (in == 126) out = -14260;
	 	 	 else if (in == 127) out = -14227;
	 	 	 else if (in == 128) out = -14195;
	 	 	 else if (in == 129) out = -14163;
	 	 	 else if (in == 130) out = -14132;
	 	 	 else if (in == 131) out = -14100;
	 	 	 else if (in == 132) out = -14069;
	 	 	 else if (in == 133) out = -14038;
	 	 	 else if (in == 134) out = -14008;
	 	 	 else if (in == 135) out = -13977;
	 	 	 else if (in == 136) out = -13947;
	 	 	 else if (in == 137) out = -13917;
	 	 	 else if (in == 138) out = -13887;
	 	 	 else if (in == 139) out = -13857;
	 	 	 else if (in == 140) out = -13828;
	 	 	 else if (in == 141) out = -13799;
	 	 	 else if (in == 142) out = -13770;
	 	 	 else if (in == 143) out = -13741;
	 	 	 else if (in == 144) out = -13713;
	 	 	 else if (in == 145) out = -13684;
	 	 	 else if (in == 146) out = -13656;
	 	 	 else if (in == 147) out = -13628;
	 	 	 else if (in == 148) out = -13600;
	 	 	 else if (in == 149) out = -13573;
	 	 	 else if (in == 150) out = -13546;
	 	 	 else if (in == 151) out = -13518;
	 	 	 else if (in == 152) out = -13491;
	 	 	 else if (in == 153) out = -13464;
	 	 	 else if (in == 154) out = -13438;
	 	 	 else if (in == 155) out = -13411;
	 	 	 else if (in == 156) out = -13385;
	 	 	 else if (in == 157) out = -13359;
	 	 	 else if (in == 158) out = -13333;
	 	 	 else if (in == 159) out = -13307;
	 	 	 else if (in == 160) out = -13281;
	 	 	 else if (in == 161) out = -13256;
	 	 	 else if (in == 162) out = -13230;
	 	 	 else if (in == 163) out = -13205;
	 	 	 else if (in == 164) out = -13180;
	 	 	 else if (in == 165) out = -13155;
	 	 	 else if (in == 166) out = -13130;
	 	 	 else if (in == 167) out = -13106;
	 	 	 else if (in == 168) out = -13081;
	 	 	 else if (in == 169) out = -13057;
	 	 	 else if (in == 170) out = -13033;
	 	 	 else if (in == 171) out = -13009;
	 	 	 else if (in == 172) out = -12985;
	 	 	 else if (in == 173) out = -12961;
	 	 	 else if (in == 174) out = -12938;
	 	 	 else if (in == 175) out = -12914;
	 	 	 else if (in == 176) out = -12891;
	 	 	 else if (in == 177) out = -12868;
	 	 	 else if (in == 178) out = -12844;
	 	 	 else if (in == 179) out = -12822;
	 	 	 else if (in == 180) out = -12799;
	 	 	 else if (in == 181) out = -12776;
	 	 	 else if (in == 182) out = -12753;
	 	 	 else if (in == 183) out = -12731;
	 	 	 else if (in == 184) out = -12709;
	 	 	 else if (in == 185) out = -12686;
	 	 	 else if (in == 186) out = -12664;
	 	 	 else if (in == 187) out = -12642;
	 	 	 else if (in == 188) out = -12621;
	 	 	 else if (in == 189) out = -12599;
	 	 	 else if (in == 190) out = -12577;
	 	 	 else if (in == 191) out = -12556;
	 	 	 else if (in == 192) out = -12534;
	 	 	 else if (in == 193) out = -12513;
	 	 	 else if (in == 194) out = -12492;
	 	 	 else if (in == 195) out = -12471;
	 	 	 else if (in == 196) out = -12450;
	 	 	 else if (in == 197) out = -12429;
	 	 	 else if (in == 198) out = -12408;
	 	 	 else if (in == 199) out = -12388;
	 	 	 else if (in == 200) out = -12367;
	 	 	 else if (in == 201) out = -12347;
	 	 	 else if (in == 202) out = -12326;
	 	 	 else if (in == 203) out = -12306;
	 	 	 else if (in == 204) out = -12286;
	 	 	 else if (in == 205) out = -12266;
	 	 	 else if (in == 206) out = -12246;
	 	 	 else if (in == 207) out = -12226;
	 	 	 else if (in == 208) out = -12207;
	 	 	 else if (in == 209) out = -12187;
	 	 	 else if (in == 210) out = -12167;
	 	 	 else if (in == 211) out = -12148;
	 	 	 else if (in == 212) out = -12128;
	 	 	 else if (in == 213) out = -12109;
	 	 	 else if (in == 214) out = -12090;
	 	 	 else if (in == 215) out = -12071;
	 	 	 else if (in == 216) out = -12052;
	 	 	 else if (in == 217) out = -12033;
	 	 	 else if (in == 218) out = -12014;
	 	 	 else if (in == 219) out = -11995;
	 	 	 else if (in == 220) out = -11977;
	 	 	 else if (in == 221) out = -11958;
	 	 	 else if (in == 222) out = -11940;
	 	 	 else if (in == 223) out = -11921;
	 	 	 else if (in == 224) out = -11903;
	 	 	 else if (in == 225) out = -11885;
	 	 	 else if (in == 226) out = -11867;
	 	 	 else if (in == 227) out = -11848;
	 	 	 else if (in == 228) out = -11830;
	 	 	 else if (in == 229) out = -11813;
	 	 	 else if (in == 230) out = -11795;
	 	 	 else if (in == 231) out = -11777;
	 	 	 else if (in == 232) out = -11759;
	 	 	 else if (in == 233) out = -11742;
	 	 	 else if (in == 234) out = -11724;
	 	 	 else if (in == 235) out = -11707;
	 	 	 else if (in == 236) out = -11689;
	 	 	 else if (in == 237) out = -11672;
	 	 	 else if (in == 238) out = -11655;
	 	 	 else if (in == 239) out = -11637;
	 	 	 else if (in == 240) out = -11620;
	 	 	 else if (in == 241) out = -11603;
	 	 	 else if (in == 242) out = -11586;
	 	 	 else if (in == 243) out = -11569;
	 	 	 else if (in == 244) out = -11553;
	 	 	 else if (in == 245) out = -11536;
	 	 	 else if (in == 246) out = -11519;
	 	 	 else if (in == 247) out = -11503;
	 	 	 else if (in == 248) out = -11486;
	 	 	 else if (in == 249) out = -11470;
	 	 	 else if (in == 250) out = -11453;
	 	 	 else if (in == 251) out = -11437;
	 	 	 else if (in == 252) out = -11421;
	 	 	 else if (in == 253) out = -11404;
	 	 	 else if (in == 254) out = -11388;
	 	 	 else if (in == 255) out = -11372;
	 	 	 else if (in == 256) out = -11356;
	 	 	 else if (in == 257) out = -11340;
	 	 	 else if (in == 258) out = -11324;
	 	 	 else if (in == 259) out = -11308;
	 	 	 else if (in == 260) out = -11293;
	 	 	 else if (in == 261) out = -11277;
	 	 	 else if (in == 262) out = -11261;
	 	 	 else if (in == 263) out = -11246;
	 	 	 else if (in == 264) out = -11230;
	 	 	 else if (in == 265) out = -11214;
	 	 	 else if (in == 266) out = -11199;
	 	 	 else if (in == 267) out = -11184;
	 	 	 else if (in == 268) out = -11168;
	 	 	 else if (in == 269) out = -11153;
	 	 	 else if (in == 270) out = -11138;
	 	 	 else if (in == 271) out = -11123;
	 	 	 else if (in == 272) out = -11108;
	 	 	 else if (in == 273) out = -11093;
	 	 	 else if (in == 274) out = -11078;
	 	 	 else if (in == 275) out = -11063;
	 	 	 else if (in == 276) out = -11048;
	 	 	 else if (in == 277) out = -11033;
	 	 	 else if (in == 278) out = -11018;
	 	 	 else if (in == 279) out = -11004;
	 	 	 else if (in == 280) out = -10989;
	 	 	 else if (in == 281) out = -10974;
	 	 	 else if (in == 282) out = -10960;
	 	 	 else if (in == 283) out = -10945;
	 	 	 else if (in == 284) out = -10931;
	 	 	 else if (in == 285) out = -10916;
	 	 	 else if (in == 286) out = -10902;
	 	 	 else if (in == 287) out = -10888;
	 	 	 else if (in == 288) out = -10874;
	 	 	 else if (in == 289) out = -10859;
	 	 	 else if (in == 290) out = -10845;
	 	 	 else if (in == 291) out = -10831;
	 	 	 else if (in == 292) out = -10817;
	 	 	 else if (in == 293) out = -10803;
	 	 	 else if (in == 294) out = -10789;
	 	 	 else if (in == 295) out = -10775;
	 	 	 else if (in == 296) out = -10761;
	 	 	 else if (in == 297) out = -10748;
	 	 	 else if (in == 298) out = -10734;
	 	 	 else if (in == 299) out = -10720;
	 	 	 else if (in == 300) out = -10706;
	 	 	 else if (in == 301) out = -10693;
	 	 	 else if (in == 302) out = -10679;
	 	 	 else if (in == 303) out = -10666;
	 	 	 else if (in == 304) out = -10652;
	 	 	 else if (in == 305) out = -10639;
	 	 	 else if (in == 306) out = -10625;
	 	 	 else if (in == 307) out = -10612;
	 	 	 else if (in == 308) out = -10599;
	 	 	 else if (in == 309) out = -10585;
	 	 	 else if (in == 310) out = -10572;
	 	 	 else if (in == 311) out = -10559;
	 	 	 else if (in == 312) out = -10546;
	 	 	 else if (in == 313) out = -10533;
	 	 	 else if (in == 314) out = -10520;
	 	 	 else if (in == 315) out = -10507;
	 	 	 else if (in == 316) out = -10494;
	 	 	 else if (in == 317) out = -10481;
	 	 	 else if (in == 318) out = -10468;
	 	 	 else if (in == 319) out = -10455;
	 	 	 else if (in == 320) out = -10442;
	 	 	 else if (in == 321) out = -10429;
	 	 	 else if (in == 322) out = -10417;
	 	 	 else if (in == 323) out = -10404;
	 	 	 else if (in == 324) out = -10391;
	 	 	 else if (in == 325) out = -10379;
	 	 	 else if (in == 326) out = -10366;
	 	 	 else if (in == 327) out = -10353;
	 	 	 else if (in == 328) out = -10341;
	 	 	 else if (in == 329) out = -10328;
	 	 	 else if (in == 330) out = -10316;
	 	 	 else if (in == 331) out = -10304;
	 	 	 else if (in == 332) out = -10291;
	 	 	 else if (in == 333) out = -10279;
	 	 	 else if (in == 334) out = -10267;
	 	 	 else if (in == 335) out = -10254;
	 	 	 else if (in == 336) out = -10242;
	 	 	 else if (in == 337) out = -10230;
	 	 	 else if (in == 338) out = -10218;
	 	 	 else if (in == 339) out = -10206;
	 	 	 else if (in == 340) out = -10194;
	 	 	 else if (in == 341) out = -10182;
	 	 	 else if (in == 342) out = -10170;
	 	 	 else if (in == 343) out = -10158;
	 	 	 else if (in == 344) out = -10146;
	 	 	 else if (in == 345) out = -10134;
	 	 	 else if (in == 346) out = -10122;
	 	 	 else if (in == 347) out = -10110;
	 	 	 else if (in == 348) out = -10098;
	 	 	 else if (in == 349) out = -10087;
	 	 	 else if (in == 350) out = -10075;
	 	 	 else if (in == 351) out = -10063;
	 	 	 else if (in == 352) out = -10052;
	 	 	 else if (in == 353) out = -10040;
	 	 	 else if (in == 354) out = -10028;
	 	 	 else if (in == 355) out = -10017;
	 	 	 else if (in == 356) out = -10005;
	 	 	 else if (in == 357) out = -9994;
	 	 	 else if (in == 358) out = -9982;
	 	 	 else if (in == 359) out = -9971;
	 	 	 else if (in == 360) out = -9960;
	 	 	 else if (in == 361) out = -9948;
	 	 	 else if (in == 362) out = -9937;
	 	 	 else if (in == 363) out = -9926;
	 	 	 else if (in == 364) out = -9914;
	 	 	 else if (in == 365) out = -9903;
	 	 	 else if (in == 366) out = -9892;
	 	 	 else if (in == 367) out = -9881;
	 	 	 else if (in == 368) out = -9870;
	 	 	 else if (in == 369) out = -9858;
	 	 	 else if (in == 370) out = -9847;
	 	 	 else if (in == 371) out = -9836;
	 	 	 else if (in == 372) out = -9825;
	 	 	 else if (in == 373) out = -9814;
	 	 	 else if (in == 374) out = -9803;
	 	 	 else if (in == 375) out = -9792;
	 	 	 else if (in == 376) out = -9781;
	 	 	 else if (in == 377) out = -9771;
	 	 	 else if (in == 378) out = -9760;
	 	 	 else if (in == 379) out = -9749;
	 	 	 else if (in == 380) out = -9738;
	 	 	 else if (in == 381) out = -9727;
	 	 	 else if (in == 382) out = -9717;
	 	 	 else if (in == 383) out = -9706;
	 	 	 else if (in == 384) out = -9695;
	 	 	 else if (in == 385) out = -9685;
	 	 	 else if (in == 386) out = -9674;
	 	 	 else if (in == 387) out = -9663;
	 	 	 else if (in == 388) out = -9653;
	 	 	 else if (in == 389) out = -9642;
	 	 	 else if (in == 390) out = -9632;
	 	 	 else if (in == 391) out = -9621;
	 	 	 else if (in == 392) out = -9611;
	 	 	 else if (in == 393) out = -9600;
	 	 	 else if (in == 394) out = -9590;
	 	 	 else if (in == 395) out = -9580;
	 	 	 else if (in == 396) out = -9569;
	 	 	 else if (in == 397) out = -9559;
	 	 	 else if (in == 398) out = -9549;
	 	 	 else if (in == 399) out = -9538;
	 	 	 else if (in == 400) out = -9528;
	 	 	 else if (in == 401) out = -9518;
	 	 	 else if (in == 402) out = -9508;
	 	 	 else if (in == 403) out = -9497;
	 	 	 else if (in == 404) out = -9487;
	 	 	 else if (in == 405) out = -9477;
	 	 	 else if (in == 406) out = -9467;
	 	 	 else if (in == 407) out = -9457;
	 	 	 else if (in == 408) out = -9447;
	 	 	 else if (in == 409) out = -9437;
	 	 	 else if (in == 410) out = -9427;
	 	 	 else if (in == 411) out = -9417;
	 	 	 else if (in == 412) out = -9407;
	 	 	 else if (in == 413) out = -9397;
	 	 	 else if (in == 414) out = -9387;
	 	 	 else if (in == 415) out = -9377;
	 	 	 else if (in == 416) out = -9367;
	 	 	 else if (in == 417) out = -9358;
	 	 	 else if (in == 418) out = -9348;
	 	 	 else if (in == 419) out = -9338;
	 	 	 else if (in == 420) out = -9328;
	 	 	 else if (in == 421) out = -9318;
	 	 	 else if (in == 422) out = -9309;
	 	 	 else if (in == 423) out = -9299;
	 	 	 else if (in == 424) out = -9289;
	 	 	 else if (in == 425) out = -9280;
	 	 	 else if (in == 426) out = -9270;
	 	 	 else if (in == 427) out = -9260;
	 	 	 else if (in == 428) out = -9251;
	 	 	 else if (in == 429) out = -9241;
	 	 	 else if (in == 430) out = -9232;
	 	 	 else if (in == 431) out = -9222;
	 	 	 else if (in == 432) out = -9213;
	 	 	 else if (in == 433) out = -9203;
	 	 	 else if (in == 434) out = -9194;
	 	 	 else if (in == 435) out = -9184;
	 	 	 else if (in == 436) out = -9175;
	 	 	 else if (in == 437) out = -9166;
	 	 	 else if (in == 438) out = -9156;
	 	 	 else if (in == 439) out = -9147;
	 	 	 else if (in == 440) out = -9138;
	 	 	 else if (in == 441) out = -9128;
	 	 	 else if (in == 442) out = -9119;
	 	 	 else if (in == 443) out = -9110;
	 	 	 else if (in == 444) out = -9101;
	 	 	 else if (in == 445) out = -9091;
	 	 	 else if (in == 446) out = -9082;
	 	 	 else if (in == 447) out = -9073;
	 	 	 else if (in == 448) out = -9064;
	 	 	 else if (in == 449) out = -9055;
	 	 	 else if (in == 450) out = -9046;
	 	 	 else if (in == 451) out = -9036;
	 	 	 else if (in == 452) out = -9027;
	 	 	 else if (in == 453) out = -9018;
	 	 	 else if (in == 454) out = -9009;
	 	 	 else if (in == 455) out = -9000;
	 	 	 else if (in == 456) out = -8991;
	 	 	 else if (in == 457) out = -8982;
	 	 	 else if (in == 458) out = -8973;
	 	 	 else if (in == 459) out = -8964;
	 	 	 else if (in == 460) out = -8956;
	 	 	 else if (in == 461) out = -8947;
	 	 	 else if (in == 462) out = -8938;
	 	 	 else if (in == 463) out = -8929;
	 	 	 else if (in == 464) out = -8920;
	 	 	 else if (in == 465) out = -8911;
	 	 	 else if (in == 466) out = -8902;
	 	 	 else if (in == 467) out = -8894;
	 	 	 else if (in == 468) out = -8885;
	 	 	 else if (in == 469) out = -8876;
	 	 	 else if (in == 470) out = -8867;
	 	 	 else if (in == 471) out = -8859;
	 	 	 else if (in == 472) out = -8850;
	 	 	 else if (in == 473) out = -8841;
	 	 	 else if (in == 474) out = -8833;
	 	 	 else if (in == 475) out = -8824;
	 	 	 else if (in == 476) out = -8816;
	 	 	 else if (in == 477) out = -8807;
	 	 	 else if (in == 478) out = -8798;
	 	 	 else if (in == 479) out = -8790;
	 	 	 else if (in == 480) out = -8781;
	 	 	 else if (in == 481) out = -8773;
	 	 	 else if (in == 482) out = -8764;
	 	 	 else if (in == 483) out = -8756;
	 	 	 else if (in == 484) out = -8747;
	 	 	 else if (in == 485) out = -8739;
	 	 	 else if (in == 486) out = -8730;
	 	 	 else if (in == 487) out = -8722;
	 	 	 else if (in == 488) out = -8714;
	 	 	 else if (in == 489) out = -8705;
	 	 	 else if (in == 490) out = -8697;
	 	 	 else if (in == 491) out = -8688;
	 	 	 else if (in == 492) out = -8680;
	 	 	 else if (in == 493) out = -8672;
	 	 	 else if (in == 494) out = -8663;
	 	 	 else if (in == 495) out = -8655;
	 	 	 else if (in == 496) out = -8647;
	 	 	 else if (in == 497) out = -8639;
	 	 	 else if (in == 498) out = -8630;
	 	 	 else if (in == 499) out = -8622;
	 	 	 else if (in == 500) out = -8614;
	 	 	 else if (in == 501) out = -8606;
	 	 	 else if (in == 502) out = -8598;
	 	 	 else if (in == 503) out = -8590;
	 	 	 else if (in == 504) out = -8581;
	 	 	 else if (in == 505) out = -8573;
	 	 	 else if (in == 506) out = -8565;
	 	 	 else if (in == 507) out = -8557;
	 	 	 else if (in == 508) out = -8549;
	 	 	 else if (in == 509) out = -8541;
	 	 	 else if (in == 510) out = -8533;
	 	 	 else if (in == 511) out = -8525;
	 	 	 else if (in == 512) out = -8517;
	 	 	 else if (in == 513) out = -8509;
	 	 	 else if (in == 514) out = -8501;
	 	 	 else if (in == 515) out = -8493;
	 	 	 else if (in == 516) out = -8485;
	 	 	 else if (in == 517) out = -8477;
	 	 	 else if (in == 518) out = -8469;
	 	 	 else if (in == 519) out = -8461;
	 	 	 else if (in == 520) out = -8453;
	 	 	 else if (in == 521) out = -8446;
	 	 	 else if (in == 522) out = -8438;
	 	 	 else if (in == 523) out = -8430;
	 	 	 else if (in == 524) out = -8422;
	 	 	 else if (in == 525) out = -8414;
	 	 	 else if (in == 526) out = -8406;
	 	 	 else if (in == 527) out = -8399;
	 	 	 else if (in == 528) out = -8391;
	 	 	 else if (in == 529) out = -8383;
	 	 	 else if (in == 530) out = -8375;
	 	 	 else if (in == 531) out = -8368;
	 	 	 else if (in == 532) out = -8360;
	 	 	 else if (in == 533) out = -8352;
	 	 	 else if (in == 534) out = -8345;
	 	 	 else if (in == 535) out = -8337;
	 	 	 else if (in == 536) out = -8329;
	 	 	 else if (in == 537) out = -8322;
	 	 	 else if (in == 538) out = -8314;
	 	 	 else if (in == 539) out = -8306;
	 	 	 else if (in == 540) out = -8299;
	 	 	 else if (in == 541) out = -8291;
	 	 	 else if (in == 542) out = -8284;
	 	 	 else if (in == 543) out = -8276;
	 	 	 else if (in == 544) out = -8269;
	 	 	 else if (in == 545) out = -8261;
	 	 	 else if (in == 546) out = -8254;
	 	 	 else if (in == 547) out = -8246;
	 	 	 else if (in == 548) out = -8239;
	 	 	 else if (in == 549) out = -8231;
	 	 	 else if (in == 550) out = -8224;
	 	 	 else if (in == 551) out = -8216;
	 	 	 else if (in == 552) out = -8209;
	 	 	 else if (in == 553) out = -8201;
	 	 	 else if (in == 554) out = -8194;
	 	 	 else if (in == 555) out = -8187;
	 	 	 else if (in == 556) out = -8179;
	 	 	 else if (in == 557) out = -8172;
	 	 	 else if (in == 558) out = -8164;
	 	 	 else if (in == 559) out = -8157;
	 	 	 else if (in == 560) out = -8150;
	 	 	 else if (in == 561) out = -8143;
	 	 	 else if (in == 562) out = -8135;
	 	 	 else if (in == 563) out = -8128;
	 	 	 else if (in == 564) out = -8121;
	 	 	 else if (in == 565) out = -8113;
	 	 	 else if (in == 566) out = -8106;
	 	 	 else if (in == 567) out = -8099;
	 	 	 else if (in == 568) out = -8092;
	 	 	 else if (in == 569) out = -8085;
	 	 	 else if (in == 570) out = -8077;
	 	 	 else if (in == 571) out = -8070;
	 	 	 else if (in == 572) out = -8063;
	 	 	 else if (in == 573) out = -8056;
	 	 	 else if (in == 574) out = -8049;
	 	 	 else if (in == 575) out = -8042;
	 	 	 else if (in == 576) out = -8034;
	 	 	 else if (in == 577) out = -8027;
	 	 	 else if (in == 578) out = -8020;
	 	 	 else if (in == 579) out = -8013;
	 	 	 else if (in == 580) out = -8006;
	 	 	 else if (in == 581) out = -7999;
	 	 	 else if (in == 582) out = -7992;
	 	 	 else if (in == 583) out = -7985;
	 	 	 else if (in == 584) out = -7978;
	 	 	 else if (in == 585) out = -7971;
	 	 	 else if (in == 586) out = -7964;
	 	 	 else if (in == 587) out = -7957;
	 	 	 else if (in == 588) out = -7950;
	 	 	 else if (in == 589) out = -7943;
	 	 	 else if (in == 590) out = -7936;
	 	 	 else if (in == 591) out = -7929;
	 	 	 else if (in == 592) out = -7922;
	 	 	 else if (in == 593) out = -7915;
	 	 	 else if (in == 594) out = -7908;
	 	 	 else if (in == 595) out = -7902;
	 	 	 else if (in == 596) out = -7895;
	 	 	 else if (in == 597) out = -7888;
	 	 	 else if (in == 598) out = -7881;
	 	 	 else if (in == 599) out = -7874;
	 	 	 else if (in == 600) out = -7867;
	 	 	 else if (in == 601) out = -7860;
	 	 	 else if (in == 602) out = -7854;
	 	 	 else if (in == 603) out = -7847;
	 	 	 else if (in == 604) out = -7840;
	 	 	 else if (in == 605) out = -7833;
	 	 	 else if (in == 606) out = -7826;
	 	 	 else if (in == 607) out = -7820;
	 	 	 else if (in == 608) out = -7813;
	 	 	 else if (in == 609) out = -7806;
	 	 	 else if (in == 610) out = -7800;
	 	 	 else if (in == 611) out = -7793;
	 	 	 else if (in == 612) out = -7786;
	 	 	 else if (in == 613) out = -7779;
	 	 	 else if (in == 614) out = -7773;
	 	 	 else if (in == 615) out = -7766;
	 	 	 else if (in == 616) out = -7759;
	 	 	 else if (in == 617) out = -7753;
	 	 	 else if (in == 618) out = -7746;
	 	 	 else if (in == 619) out = -7740;
	 	 	 else if (in == 620) out = -7733;
	 	 	 else if (in == 621) out = -7726;
	 	 	 else if (in == 622) out = -7720;
	 	 	 else if (in == 623) out = -7713;
	 	 	 else if (in == 624) out = -7707;
	 	 	 else if (in == 625) out = -7700;
	 	 	 else if (in == 626) out = -7693;
	 	 	 else if (in == 627) out = -7687;
	 	 	 else if (in == 628) out = -7680;
	 	 	 else if (in == 629) out = -7674;
	 	 	 else if (in == 630) out = -7667;
	 	 	 else if (in == 631) out = -7661;
	 	 	 else if (in == 632) out = -7654;
	 	 	 else if (in == 633) out = -7648;
	 	 	 else if (in == 634) out = -7641;
	 	 	 else if (in == 635) out = -7635;
	 	 	 else if (in == 636) out = -7629;
	 	 	 else if (in == 637) out = -7622;
	 	 	 else if (in == 638) out = -7616;
	 	 	 else if (in == 639) out = -7609;
	 	 	 else if (in == 640) out = -7603;
	 	 	 else if (in == 641) out = -7597;
	 	 	 else if (in == 642) out = -7590;
	 	 	 else if (in == 643) out = -7584;
	 	 	 else if (in == 644) out = -7577;
	 	 	 else if (in == 645) out = -7571;
	 	 	 else if (in == 646) out = -7565;
	 	 	 else if (in == 647) out = -7558;
	 	 	 else if (in == 648) out = -7552;
	 	 	 else if (in == 649) out = -7546;
	 	 	 else if (in == 650) out = -7539;
	 	 	 else if (in == 651) out = -7533;
	 	 	 else if (in == 652) out = -7527;
	 	 	 else if (in == 653) out = -7521;
	 	 	 else if (in == 654) out = -7514;
	 	 	 else if (in == 655) out = -7508;
	 	 	 else if (in == 656) out = -7502;
	 	 	 else if (in == 657) out = -7496;
	 	 	 else if (in == 658) out = -7489;
	 	 	 else if (in == 659) out = -7483;
	 	 	 else if (in == 660) out = -7477;
	 	 	 else if (in == 661) out = -7471;
	 	 	 else if (in == 662) out = -7464;
	 	 	 else if (in == 663) out = -7458;
	 	 	 else if (in == 664) out = -7452;
	 	 	 else if (in == 665) out = -7446;
	 	 	 else if (in == 666) out = -7440;
	 	 	 else if (in == 667) out = -7434;
	 	 	 else if (in == 668) out = -7428;
	 	 	 else if (in == 669) out = -7421;
	 	 	 else if (in == 670) out = -7415;
	 	 	 else if (in == 671) out = -7409;
	 	 	 else if (in == 672) out = -7403;
	 	 	 else if (in == 673) out = -7397;
	 	 	 else if (in == 674) out = -7391;
	 	 	 else if (in == 675) out = -7385;
	 	 	 else if (in == 676) out = -7379;
	 	 	 else if (in == 677) out = -7373;
	 	 	 else if (in == 678) out = -7367;
	 	 	 else if (in == 679) out = -7361;
	 	 	 else if (in == 680) out = -7355;
	 	 	 else if (in == 681) out = -7349;
	 	 	 else if (in == 682) out = -7343;
	 	 	 else if (in == 683) out = -7337;
	 	 	 else if (in == 684) out = -7331;
	 	 	 else if (in == 685) out = -7325;
	 	 	 else if (in == 686) out = -7319;
	 	 	 else if (in == 687) out = -7313;
	 	 	 else if (in == 688) out = -7307;
	 	 	 else if (in == 689) out = -7301;
	 	 	 else if (in == 690) out = -7295;
	 	 	 else if (in == 691) out = -7289;
	 	 	 else if (in == 692) out = -7283;
	 	 	 else if (in == 693) out = -7277;
	 	 	 else if (in == 694) out = -7271;
	 	 	 else if (in == 695) out = -7265;
	 	 	 else if (in == 696) out = -7259;
	 	 	 else if (in == 697) out = -7253;
	 	 	 else if (in == 698) out = -7248;
	 	 	 else if (in == 699) out = -7242;
	 	 	 else if (in == 700) out = -7236;
	 	 	 else if (in == 701) out = -7230;
	 	 	 else if (in == 702) out = -7224;
	 	 	 else if (in == 703) out = -7218;
	 	 	 else if (in == 704) out = -7213;
	 	 	 else if (in == 705) out = -7207;
	 	 	 else if (in == 706) out = -7201;
	 	 	 else if (in == 707) out = -7195;
	 	 	 else if (in == 708) out = -7189;
	 	 	 else if (in == 709) out = -7184;
	 	 	 else if (in == 710) out = -7178;
	 	 	 else if (in == 711) out = -7172;
	 	 	 else if (in == 712) out = -7166;
	 	 	 else if (in == 713) out = -7160;
	 	 	 else if (in == 714) out = -7155;
	 	 	 else if (in == 715) out = -7149;
	 	 	 else if (in == 716) out = -7143;
	 	 	 else if (in == 717) out = -7138;
	 	 	 else if (in == 718) out = -7132;
	 	 	 else if (in == 719) out = -7126;
	 	 	 else if (in == 720) out = -7120;
	 	 	 else if (in == 721) out = -7115;
	 	 	 else if (in == 722) out = -7109;
	 	 	 else if (in == 723) out = -7103;
	 	 	 else if (in == 724) out = -7098;
	 	 	 else if (in == 725) out = -7092;
	 	 	 else if (in == 726) out = -7086;
	 	 	 else if (in == 727) out = -7081;
	 	 	 else if (in == 728) out = -7075;
	 	 	 else if (in == 729) out = -7070;
	 	 	 else if (in == 730) out = -7064;
	 	 	 else if (in == 731) out = -7058;
	 	 	 else if (in == 732) out = -7053;
	 	 	 else if (in == 733) out = -7047;
	 	 	 else if (in == 734) out = -7042;
	 	 	 else if (in == 735) out = -7036;
	 	 	 else if (in == 736) out = -7030;
	 	 	 else if (in == 737) out = -7025;
	 	 	 else if (in == 738) out = -7019;
	 	 	 else if (in == 739) out = -7014;
	 	 	 else if (in == 740) out = -7008;
	 	 	 else if (in == 741) out = -7003;
	 	 	 else if (in == 742) out = -6997;
	 	 	 else if (in == 743) out = -6992;
	 	 	 else if (in == 744) out = -6986;
	 	 	 else if (in == 745) out = -6981;
	 	 	 else if (in == 746) out = -6975;
	 	 	 else if (in == 747) out = -6970;
	 	 	 else if (in == 748) out = -6964;
	 	 	 else if (in == 749) out = -6959;
	 	 	 else if (in == 750) out = -6953;
	 	 	 else if (in == 751) out = -6948;
	 	 	 else if (in == 752) out = -6942;
	 	 	 else if (in == 753) out = -6937;
	 	 	 else if (in == 754) out = -6931;
	 	 	 else if (in == 755) out = -6926;
	 	 	 else if (in == 756) out = -6921;
	 	 	 else if (in == 757) out = -6915;
	 	 	 else if (in == 758) out = -6910;
	 	 	 else if (in == 759) out = -6904;
	 	 	 else if (in == 760) out = -6899;
	 	 	 else if (in == 761) out = -6894;
	 	 	 else if (in == 762) out = -6888;
	 	 	 else if (in == 763) out = -6883;
	 	 	 else if (in == 764) out = -6877;
	 	 	 else if (in == 765) out = -6872;
	 	 	 else if (in == 766) out = -6867;
	 	 	 else if (in == 767) out = -6861;
	 	 	 else if (in == 768) out = -6856;
	 	 	 else if (in == 769) out = -6851;
	 	 	 else if (in == 770) out = -6845;
	 	 	 else if (in == 771) out = -6840;
	 	 	 else if (in == 772) out = -6835;
	 	 	 else if (in == 773) out = -6830;
	 	 	 else if (in == 774) out = -6824;
	 	 	 else if (in == 775) out = -6819;
	 	 	 else if (in == 776) out = -6814;
	 	 	 else if (in == 777) out = -6808;
	 	 	 else if (in == 778) out = -6803;
	 	 	 else if (in == 779) out = -6798;
	 	 	 else if (in == 780) out = -6793;
	 	 	 else if (in == 781) out = -6787;
	 	 	 else if (in == 782) out = -6782;
	 	 	 else if (in == 783) out = -6777;
	 	 	 else if (in == 784) out = -6772;
	 	 	 else if (in == 785) out = -6766;
	 	 	 else if (in == 786) out = -6761;
	 	 	 else if (in == 787) out = -6756;
	 	 	 else if (in == 788) out = -6751;
	 	 	 else if (in == 789) out = -6746;
	 	 	 else if (in == 790) out = -6740;
	 	 	 else if (in == 791) out = -6735;
	 	 	 else if (in == 792) out = -6730;
	 	 	 else if (in == 793) out = -6725;
	 	 	 else if (in == 794) out = -6720;
	 	 	 else if (in == 795) out = -6715;
	 	 	 else if (in == 796) out = -6709;
	 	 	 else if (in == 797) out = -6704;
	 	 	 else if (in == 798) out = -6699;
	 	 	 else if (in == 799) out = -6694;
	 	 	 else if (in == 800) out = -6689;
	 	 	 else if (in == 801) out = -6684;
	 	 	 else if (in == 802) out = -6679;
	 	 	 else if (in == 803) out = -6674;
	 	 	 else if (in == 804) out = -6668;
	 	 	 else if (in == 805) out = -6663;
	 	 	 else if (in == 806) out = -6658;
	 	 	 else if (in == 807) out = -6653;
	 	 	 else if (in == 808) out = -6648;
	 	 	 else if (in == 809) out = -6643;
	 	 	 else if (in == 810) out = -6638;
	 	 	 else if (in == 811) out = -6633;
	 	 	 else if (in == 812) out = -6628;
	 	 	 else if (in == 813) out = -6623;
	 	 	 else if (in == 814) out = -6618;
	 	 	 else if (in == 815) out = -6613;
	 	 	 else if (in == 816) out = -6608;
	 	 	 else if (in == 817) out = -6603;
	 	 	 else if (in == 818) out = -6598;
	 	 	 else if (in == 819) out = -6593;
	 	 	 else if (in == 820) out = -6588;
	 	 	 else if (in == 821) out = -6583;
	 	 	 else if (in == 822) out = -6578;
	 	 	 else if (in == 823) out = -6573;
	 	 	 else if (in == 824) out = -6568;
	 	 	 else if (in == 825) out = -6563;
	 	 	 else if (in == 826) out = -6558;
	 	 	 else if (in == 827) out = -6553;
	 	 	 else if (in == 828) out = -6548;
	 	 	 else if (in == 829) out = -6543;
	 	 	 else if (in == 830) out = -6538;
	 	 	 else if (in == 831) out = -6533;
	 	 	 else if (in == 832) out = -6528;
	 	 	 else if (in == 833) out = -6523;
	 	 	 else if (in == 834) out = -6518;
	 	 	 else if (in == 835) out = -6514;
	 	 	 else if (in == 836) out = -6509;
	 	 	 else if (in == 837) out = -6504;
	 	 	 else if (in == 838) out = -6499;
	 	 	 else if (in == 839) out = -6494;
	 	 	 else if (in == 840) out = -6489;
	 	 	 else if (in == 841) out = -6484;
	 	 	 else if (in == 842) out = -6479;
	 	 	 else if (in == 843) out = -6474;
	 	 	 else if (in == 844) out = -6470;
	 	 	 else if (in == 845) out = -6465;
	 	 	 else if (in == 846) out = -6460;
	 	 	 else if (in == 847) out = -6455;
	 	 	 else if (in == 848) out = -6450;
	 	 	 else if (in == 849) out = -6445;
	 	 	 else if (in == 850) out = -6441;
	 	 	 else if (in == 851) out = -6436;
	 	 	 else if (in == 852) out = -6431;
	 	 	 else if (in == 853) out = -6426;
	 	 	 else if (in == 854) out = -6421;
	 	 	 else if (in == 855) out = -6417;
	 	 	 else if (in == 856) out = -6412;
	 	 	 else if (in == 857) out = -6407;
	 	 	 else if (in == 858) out = -6402;
	 	 	 else if (in == 859) out = -6397;
	 	 	 else if (in == 860) out = -6393;
	 	 	 else if (in == 861) out = -6388;
	 	 	 else if (in == 862) out = -6383;
	 	 	 else if (in == 863) out = -6378;
	 	 	 else if (in == 864) out = -6374;
	 	 	 else if (in == 865) out = -6369;
	 	 	 else if (in == 866) out = -6364;
	 	 	 else if (in == 867) out = -6359;
	 	 	 else if (in == 868) out = -6355;
	 	 	 else if (in == 869) out = -6350;
	 	 	 else if (in == 870) out = -6345;
	 	 	 else if (in == 871) out = -6341;
	 	 	 else if (in == 872) out = -6336;
	 	 	 else if (in == 873) out = -6331;
	 	 	 else if (in == 874) out = -6327;
	 	 	 else if (in == 875) out = -6322;
	 	 	 else if (in == 876) out = -6317;
	 	 	 else if (in == 877) out = -6312;
	 	 	 else if (in == 878) out = -6308;
	 	 	 else if (in == 879) out = -6303;
	 	 	 else if (in == 880) out = -6299;
	 	 	 else if (in == 881) out = -6294;
	 	 	 else if (in == 882) out = -6289;
	 	 	 else if (in == 883) out = -6285;
	 	 	 else if (in == 884) out = -6280;
	 	 	 else if (in == 885) out = -6275;
	 	 	 else if (in == 886) out = -6271;
	 	 	 else if (in == 887) out = -6266;
	 	 	 else if (in == 888) out = -6261;
	 	 	 else if (in == 889) out = -6257;
	 	 	 else if (in == 890) out = -6252;
	 	 	 else if (in == 891) out = -6248;
	 	 	 else if (in == 892) out = -6243;
	 	 	 else if (in == 893) out = -6238;
	 	 	 else if (in == 894) out = -6234;
	 	 	 else if (in == 895) out = -6229;
	 	 	 else if (in == 896) out = -6225;
	 	 	 else if (in == 897) out = -6220;
	 	 	 else if (in == 898) out = -6216;
	 	 	 else if (in == 899) out = -6211;
	 	 	 else if (in == 900) out = -6206;
	 	 	 else if (in == 901) out = -6202;
	 	 	 else if (in == 902) out = -6197;
	 	 	 else if (in == 903) out = -6193;
	 	 	 else if (in == 904) out = -6188;
	 	 	 else if (in == 905) out = -6184;
	 	 	 else if (in == 906) out = -6179;
	 	 	 else if (in == 907) out = -6175;
	 	 	 else if (in == 908) out = -6170;
	 	 	 else if (in == 909) out = -6166;
	 	 	 else if (in == 910) out = -6161;
	 	 	 else if (in == 911) out = -6157;
	 	 	 else if (in == 912) out = -6152;
	 	 	 else if (in == 913) out = -6148;
	 	 	 else if (in == 914) out = -6143;
	 	 	 else if (in == 915) out = -6139;
	 	 	 else if (in == 916) out = -6134;
	 	 	 else if (in == 917) out = -6130;
	 	 	 else if (in == 918) out = -6125;
	 	 	 else if (in == 919) out = -6121;
	 	 	 else if (in == 920) out = -6116;
	 	 	 else if (in == 921) out = -6112;
	 	 	 else if (in == 922) out = -6108;
	 	 	 else if (in == 923) out = -6103;
	 	 	 else if (in == 924) out = -6099;
	 	 	 else if (in == 925) out = -6094;
	 	 	 else if (in == 926) out = -6090;
	 	 	 else if (in == 927) out = -6085;
	 	 	 else if (in == 928) out = -6081;
	 	 	 else if (in == 929) out = -6077;
	 	 	 else if (in == 930) out = -6072;
	 	 	 else if (in == 931) out = -6068;
	 	 	 else if (in == 932) out = -6063;
	 	 	 else if (in == 933) out = -6059;
	 	 	 else if (in == 934) out = -6055;
	 	 	 else if (in == 935) out = -6050;
	 	 	 else if (in == 936) out = -6046;
	 	 	 else if (in == 937) out = -6041;
	 	 	 else if (in == 938) out = -6037;
	 	 	 else if (in == 939) out = -6033;
	 	 	 else if (in == 940) out = -6028;
	 	 	 else if (in == 941) out = -6024;
	 	 	 else if (in == 942) out = -6020;
	 	 	 else if (in == 943) out = -6015;
	 	 	 else if (in == 944) out = -6011;
	 	 	 else if (in == 945) out = -6007;
	 	 	 else if (in == 946) out = -6002;
	 	 	 else if (in == 947) out = -5998;
	 	 	 else if (in == 948) out = -5994;
	 	 	 else if (in == 949) out = -5989;
	 	 	 else if (in == 950) out = -5985;
	 	 	 else if (in == 951) out = -5981;
	 	 	 else if (in == 952) out = -5976;
	 	 	 else if (in == 953) out = -5972;
	 	 	 else if (in == 954) out = -5968;
	 	 	 else if (in == 955) out = -5964;
	 	 	 else if (in == 956) out = -5959;
	 	 	 else if (in == 957) out = -5955;
	 	 	 else if (in == 958) out = -5951;
	 	 	 else if (in == 959) out = -5946;
	 	 	 else if (in == 960) out = -5942;
	 	 	 else if (in == 961) out = -5938;
	 	 	 else if (in == 962) out = -5934;
	 	 	 else if (in == 963) out = -5929;
	 	 	 else if (in == 964) out = -5925;
	 	 	 else if (in == 965) out = -5921;
	 	 	 else if (in == 966) out = -5917;
	 	 	 else if (in == 967) out = -5912;
	 	 	 else if (in == 968) out = -5908;
	 	 	 else if (in == 969) out = -5904;
	 	 	 else if (in == 970) out = -5900;
	 	 	 else if (in == 971) out = -5895;
	 	 	 else if (in == 972) out = -5891;
	 	 	 else if (in == 973) out = -5887;
	 	 	 else if (in == 974) out = -5883;
	 	 	 else if (in == 975) out = -5879;
	 	 	 else if (in == 976) out = -5874;
	 	 	 else if (in == 977) out = -5870;
	 	 	 else if (in == 978) out = -5866;
	 	 	 else if (in == 979) out = -5862;
	 	 	 else if (in == 980) out = -5858;
	 	 	 else if (in == 981) out = -5853;
	 	 	 else if (in == 982) out = -5849;
	 	 	 else if (in == 983) out = -5845;
	 	 	 else if (in == 984) out = -5841;
	 	 	 else if (in == 985) out = -5837;
	 	 	 else if (in == 986) out = -5833;
	 	 	 else if (in == 987) out = -5829;
	 	 	 else if (in == 988) out = -5824;
	 	 	 else if (in == 989) out = -5820;
	 	 	 else if (in == 990) out = -5816;
	 	 	 else if (in == 991) out = -5812;
	 	 	 else if (in == 992) out = -5808;
	 	 	 else if (in == 993) out = -5804;
	 	 	 else if (in == 994) out = -5800;
	 	 	 else if (in == 995) out = -5795;
	 	 	 else if (in == 996) out = -5791;
	 	 	 else if (in == 997) out = -5787;
	 	 	 else if (in == 998) out = -5783;
	 	 	 else if (in == 999) out = -5779;
	 	 	 else if (in == 1000) out = -5775;
	 	 	 else if (in == 1001) out = -5771;
	 	 	 else if (in == 1002) out = -5767;
	 	 	 else if (in == 1003) out = -5763;
	 	 	 else if (in == 1004) out = -5759;
	 	 	 else if (in == 1005) out = -5754;
	 	 	 else if (in == 1006) out = -5750;
	 	 	 else if (in == 1007) out = -5746;
	 	 	 else if (in == 1008) out = -5742;
	 	 	 else if (in == 1009) out = -5738;
	 	 	 else if (in == 1010) out = -5734;
	 	 	 else if (in == 1011) out = -5730;
	 	 	 else if (in == 1012) out = -5726;
	 	 	 else if (in == 1013) out = -5722;
	 	 	 else if (in == 1014) out = -5718;
	 	 	 else if (in == 1015) out = -5714;
	 	 	 else if (in == 1016) out = -5710;
	 	 	 else if (in == 1017) out = -5706;
	 	 	 else if (in == 1018) out = -5702;
	 	 	 else if (in == 1019) out = -5698;
	 	 	 else if (in == 1020) out = -5694;
	 	 	 else if (in == 1021) out = -5690;
	 	 	 else if (in == 1022) out = -5686;
	 	 	 else if (in == 1023) out = -5682;
	 	 	 else if (in == 1024) out = -5678;
	 	 	 else if (in == 1025) out = -5674;
	 	 	 else if (in == 1026) out = -5670;
	 	 	 else if (in == 1027) out = -5666;
	 	 	 else if (in == 1028) out = -5662;
	 	 	 else if (in == 1029) out = -5658;
	 	 	 else if (in == 1030) out = -5654;
	 	 	 else if (in == 1031) out = -5650;
	 	 	 else if (in == 1032) out = -5646;
	 	 	 else if (in == 1033) out = -5642;
	 	 	 else if (in == 1034) out = -5638;
	 	 	 else if (in == 1035) out = -5634;
	 	 	 else if (in == 1036) out = -5630;
	 	 	 else if (in == 1037) out = -5626;
	 	 	 else if (in == 1038) out = -5622;
	 	 	 else if (in == 1039) out = -5618;
	 	 	 else if (in == 1040) out = -5614;
	 	 	 else if (in == 1041) out = -5610;
	 	 	 else if (in == 1042) out = -5606;
	 	 	 else if (in == 1043) out = -5602;
	 	 	 else if (in == 1044) out = -5599;
	 	 	 else if (in == 1045) out = -5595;
	 	 	 else if (in == 1046) out = -5591;
	 	 	 else if (in == 1047) out = -5587;
	 	 	 else if (in == 1048) out = -5583;
	 	 	 else if (in == 1049) out = -5579;
	 	 	 else if (in == 1050) out = -5575;
	 	 	 else if (in == 1051) out = -5571;
	 	 	 else if (in == 1052) out = -5567;
	 	 	 else if (in == 1053) out = -5563;
	 	 	 else if (in == 1054) out = -5559;
	 	 	 else if (in == 1055) out = -5556;
	 	 	 else if (in == 1056) out = -5552;
	 	 	 else if (in == 1057) out = -5548;
	 	 	 else if (in == 1058) out = -5544;
	 	 	 else if (in == 1059) out = -5540;
	 	 	 else if (in == 1060) out = -5536;
	 	 	 else if (in == 1061) out = -5532;
	 	 	 else if (in == 1062) out = -5529;
	 	 	 else if (in == 1063) out = -5525;
	 	 	 else if (in == 1064) out = -5521;
	 	 	 else if (in == 1065) out = -5517;
	 	 	 else if (in == 1066) out = -5513;
	 	 	 else if (in == 1067) out = -5509;
	 	 	 else if (in == 1068) out = -5505;
	 	 	 else if (in == 1069) out = -5502;
	 	 	 else if (in == 1070) out = -5498;
	 	 	 else if (in == 1071) out = -5494;
	 	 	 else if (in == 1072) out = -5490;
	 	 	 else if (in == 1073) out = -5486;
	 	 	 else if (in == 1074) out = -5482;
	 	 	 else if (in == 1075) out = -5479;
	 	 	 else if (in == 1076) out = -5475;
	 	 	 else if (in == 1077) out = -5471;
	 	 	 else if (in == 1078) out = -5467;
	 	 	 else if (in == 1079) out = -5463;
	 	 	 else if (in == 1080) out = -5460;
	 	 	 else if (in == 1081) out = -5456;
	 	 	 else if (in == 1082) out = -5452;
	 	 	 else if (in == 1083) out = -5448;
	 	 	 else if (in == 1084) out = -5445;
	 	 	 else if (in == 1085) out = -5441;
	 	 	 else if (in == 1086) out = -5437;
	 	 	 else if (in == 1087) out = -5433;
	 	 	 else if (in == 1088) out = -5429;
	 	 	 else if (in == 1089) out = -5426;
	 	 	 else if (in == 1090) out = -5422;
	 	 	 else if (in == 1091) out = -5418;
	 	 	 else if (in == 1092) out = -5414;
	 	 	 else if (in == 1093) out = -5411;
	 	 	 else if (in == 1094) out = -5407;
	 	 	 else if (in == 1095) out = -5403;
	 	 	 else if (in == 1096) out = -5399;
	 	 	 else if (in == 1097) out = -5396;
	 	 	 else if (in == 1098) out = -5392;
	 	 	 else if (in == 1099) out = -5388;
	 	 	 else if (in == 1100) out = -5385;
	 	 	 else if (in == 1101) out = -5381;
	 	 	 else if (in == 1102) out = -5377;
	 	 	 else if (in == 1103) out = -5373;
	 	 	 else if (in == 1104) out = -5370;
	 	 	 else if (in == 1105) out = -5366;
	 	 	 else if (in == 1106) out = -5362;
	 	 	 else if (in == 1107) out = -5359;
	 	 	 else if (in == 1108) out = -5355;
	 	 	 else if (in == 1109) out = -5351;
	 	 	 else if (in == 1110) out = -5347;
	 	 	 else if (in == 1111) out = -5344;
	 	 	 else if (in == 1112) out = -5340;
	 	 	 else if (in == 1113) out = -5336;
	 	 	 else if (in == 1114) out = -5333;
	 	 	 else if (in == 1115) out = -5329;
	 	 	 else if (in == 1116) out = -5325;
	 	 	 else if (in == 1117) out = -5322;
	 	 	 else if (in == 1118) out = -5318;
	 	 	 else if (in == 1119) out = -5314;
	 	 	 else if (in == 1120) out = -5311;
	 	 	 else if (in == 1121) out = -5307;
	 	 	 else if (in == 1122) out = -5303;
	 	 	 else if (in == 1123) out = -5300;
	 	 	 else if (in == 1124) out = -5296;
	 	 	 else if (in == 1125) out = -5292;
	 	 	 else if (in == 1126) out = -5289;
	 	 	 else if (in == 1127) out = -5285;
	 	 	 else if (in == 1128) out = -5282;
	 	 	 else if (in == 1129) out = -5278;
	 	 	 else if (in == 1130) out = -5274;
	 	 	 else if (in == 1131) out = -5271;
	 	 	 else if (in == 1132) out = -5267;
	 	 	 else if (in == 1133) out = -5263;
	 	 	 else if (in == 1134) out = -5260;
	 	 	 else if (in == 1135) out = -5256;
	 	 	 else if (in == 1136) out = -5253;
	 	 	 else if (in == 1137) out = -5249;
	 	 	 else if (in == 1138) out = -5245;
	 	 	 else if (in == 1139) out = -5242;
	 	 	 else if (in == 1140) out = -5238;
	 	 	 else if (in == 1141) out = -5235;
	 	 	 else if (in == 1142) out = -5231;
	 	 	 else if (in == 1143) out = -5227;
	 	 	 else if (in == 1144) out = -5224;
	 	 	 else if (in == 1145) out = -5220;
	 	 	 else if (in == 1146) out = -5217;
	 	 	 else if (in == 1147) out = -5213;
	 	 	 else if (in == 1148) out = -5210;
	 	 	 else if (in == 1149) out = -5206;
	 	 	 else if (in == 1150) out = -5202;
	 	 	 else if (in == 1151) out = -5199;
	 	 	 else if (in == 1152) out = -5195;
	 	 	 else if (in == 1153) out = -5192;
	 	 	 else if (in == 1154) out = -5188;
	 	 	 else if (in == 1155) out = -5185;
	 	 	 else if (in == 1156) out = -5181;
	 	 	 else if (in == 1157) out = -5178;
	 	 	 else if (in == 1158) out = -5174;
	 	 	 else if (in == 1159) out = -5171;
	 	 	 else if (in == 1160) out = -5167;
	 	 	 else if (in == 1161) out = -5163;
	 	 	 else if (in == 1162) out = -5160;
	 	 	 else if (in == 1163) out = -5156;
	 	 	 else if (in == 1164) out = -5153;
	 	 	 else if (in == 1165) out = -5149;
	 	 	 else if (in == 1166) out = -5146;
	 	 	 else if (in == 1167) out = -5142;
	 	 	 else if (in == 1168) out = -5139;
	 	 	 else if (in == 1169) out = -5135;
	 	 	 else if (in == 1170) out = -5132;
	 	 	 else if (in == 1171) out = -5128;
	 	 	 else if (in == 1172) out = -5125;
	 	 	 else if (in == 1173) out = -5121;
	 	 	 else if (in == 1174) out = -5118;
	 	 	 else if (in == 1175) out = -5114;
	 	 	 else if (in == 1176) out = -5111;
	 	 	 else if (in == 1177) out = -5107;
	 	 	 else if (in == 1178) out = -5104;
	 	 	 else if (in == 1179) out = -5100;
	 	 	 else if (in == 1180) out = -5097;
	 	 	 else if (in == 1181) out = -5093;
	 	 	 else if (in == 1182) out = -5090;
	 	 	 else if (in == 1183) out = -5087;
	 	 	 else if (in == 1184) out = -5083;
	 	 	 else if (in == 1185) out = -5080;
	 	 	 else if (in == 1186) out = -5076;
	 	 	 else if (in == 1187) out = -5073;
	 	 	 else if (in == 1188) out = -5069;
	 	 	 else if (in == 1189) out = -5066;
	 	 	 else if (in == 1190) out = -5062;
	 	 	 else if (in == 1191) out = -5059;
	 	 	 else if (in == 1192) out = -5056;
	 	 	 else if (in == 1193) out = -5052;
	 	 	 else if (in == 1194) out = -5049;
	 	 	 else if (in == 1195) out = -5045;
	 	 	 else if (in == 1196) out = -5042;
	 	 	 else if (in == 1197) out = -5038;
	 	 	 else if (in == 1198) out = -5035;
	 	 	 else if (in == 1199) out = -5032;
	 	 	 else if (in == 1200) out = -5028;
	 	 	 else if (in == 1201) out = -5025;
	 	 	 else if (in == 1202) out = -5021;
	 	 	 else if (in == 1203) out = -5018;
	 	 	 else if (in == 1204) out = -5014;
	 	 	 else if (in == 1205) out = -5011;
	 	 	 else if (in == 1206) out = -5008;
	 	 	 else if (in == 1207) out = -5004;
	 	 	 else if (in == 1208) out = -5001;
	 	 	 else if (in == 1209) out = -4998;
	 	 	 else if (in == 1210) out = -4994;
	 	 	 else if (in == 1211) out = -4991;
	 	 	 else if (in == 1212) out = -4987;
	 	 	 else if (in == 1213) out = -4984;
	 	 	 else if (in == 1214) out = -4981;
	 	 	 else if (in == 1215) out = -4977;
	 	 	 else if (in == 1216) out = -4974;
	 	 	 else if (in == 1217) out = -4970;
	 	 	 else if (in == 1218) out = -4967;
	 	 	 else if (in == 1219) out = -4964;
	 	 	 else if (in == 1220) out = -4960;
	 	 	 else if (in == 1221) out = -4957;
	 	 	 else if (in == 1222) out = -4954;
	 	 	 else if (in == 1223) out = -4950;
	 	 	 else if (in == 1224) out = -4947;
	 	 	 else if (in == 1225) out = -4944;
	 	 	 else if (in == 1226) out = -4940;
	 	 	 else if (in == 1227) out = -4937;
	 	 	 else if (in == 1228) out = -4934;
	 	 	 else if (in == 1229) out = -4930;
	 	 	 else if (in == 1230) out = -4927;
	 	 	 else if (in == 1231) out = -4924;
	 	 	 else if (in == 1232) out = -4920;
	 	 	 else if (in == 1233) out = -4917;
	 	 	 else if (in == 1234) out = -4914;
	 	 	 else if (in == 1235) out = -4910;
	 	 	 else if (in == 1236) out = -4907;
	 	 	 else if (in == 1237) out = -4904;
	 	 	 else if (in == 1238) out = -4900;
	 	 	 else if (in == 1239) out = -4897;
	 	 	 else if (in == 1240) out = -4894;
	 	 	 else if (in == 1241) out = -4891;
	 	 	 else if (in == 1242) out = -4887;
	 	 	 else if (in == 1243) out = -4884;
	 	 	 else if (in == 1244) out = -4881;
	 	 	 else if (in == 1245) out = -4877;
	 	 	 else if (in == 1246) out = -4874;
	 	 	 else if (in == 1247) out = -4871;
	 	 	 else if (in == 1248) out = -4867;
	 	 	 else if (in == 1249) out = -4864;
	 	 	 else if (in == 1250) out = -4861;
	 	 	 else if (in == 1251) out = -4858;
	 	 	 else if (in == 1252) out = -4854;
	 	 	 else if (in == 1253) out = -4851;
	 	 	 else if (in == 1254) out = -4848;
	 	 	 else if (in == 1255) out = -4845;
	 	 	 else if (in == 1256) out = -4841;
	 	 	 else if (in == 1257) out = -4838;
	 	 	 else if (in == 1258) out = -4835;
	 	 	 else if (in == 1259) out = -4832;
	 	 	 else if (in == 1260) out = -4828;
	 	 	 else if (in == 1261) out = -4825;
	 	 	 else if (in == 1262) out = -4822;
	 	 	 else if (in == 1263) out = -4819;
	 	 	 else if (in == 1264) out = -4815;
	 	 	 else if (in == 1265) out = -4812;
	 	 	 else if (in == 1266) out = -4809;
	 	 	 else if (in == 1267) out = -4806;
	 	 	 else if (in == 1268) out = -4802;
	 	 	 else if (in == 1269) out = -4799;
	 	 	 else if (in == 1270) out = -4796;
	 	 	 else if (in == 1271) out = -4793;
	 	 	 else if (in == 1272) out = -4789;
	 	 	 else if (in == 1273) out = -4786;
	 	 	 else if (in == 1274) out = -4783;
	 	 	 else if (in == 1275) out = -4780;
	 	 	 else if (in == 1276) out = -4777;
	 	 	 else if (in == 1277) out = -4773;
	 	 	 else if (in == 1278) out = -4770;
	 	 	 else if (in == 1279) out = -4767;
	 	 	 else if (in == 1280) out = -4764;
	 	 	 else if (in == 1281) out = -4761;
	 	 	 else if (in == 1282) out = -4757;
	 	 	 else if (in == 1283) out = -4754;
	 	 	 else if (in == 1284) out = -4751;
	 	 	 else if (in == 1285) out = -4748;
	 	 	 else if (in == 1286) out = -4745;
	 	 	 else if (in == 1287) out = -4741;
	 	 	 else if (in == 1288) out = -4738;
	 	 	 else if (in == 1289) out = -4735;
	 	 	 else if (in == 1290) out = -4732;
	 	 	 else if (in == 1291) out = -4729;
	 	 	 else if (in == 1292) out = -4726;
	 	 	 else if (in == 1293) out = -4722;
	 	 	 else if (in == 1294) out = -4719;
	 	 	 else if (in == 1295) out = -4716;
	 	 	 else if (in == 1296) out = -4713;
	 	 	 else if (in == 1297) out = -4710;
	 	 	 else if (in == 1298) out = -4707;
	 	 	 else if (in == 1299) out = -4703;
	 	 	 else if (in == 1300) out = -4700;
	 	 	 else if (in == 1301) out = -4697;
	 	 	 else if (in == 1302) out = -4694;
	 	 	 else if (in == 1303) out = -4691;
	 	 	 else if (in == 1304) out = -4688;
	 	 	 else if (in == 1305) out = -4685;
	 	 	 else if (in == 1306) out = -4681;
	 	 	 else if (in == 1307) out = -4678;
	 	 	 else if (in == 1308) out = -4675;
	 	 	 else if (in == 1309) out = -4672;
	 	 	 else if (in == 1310) out = -4669;
	 	 	 else if (in == 1311) out = -4666;
	 	 	 else if (in == 1312) out = -4663;
	 	 	 else if (in == 1313) out = -4660;
	 	 	 else if (in == 1314) out = -4656;
	 	 	 else if (in == 1315) out = -4653;
	 	 	 else if (in == 1316) out = -4650;
	 	 	 else if (in == 1317) out = -4647;
	 	 	 else if (in == 1318) out = -4644;
	 	 	 else if (in == 1319) out = -4641;
	 	 	 else if (in == 1320) out = -4638;
	 	 	 else if (in == 1321) out = -4635;
	 	 	 else if (in == 1322) out = -4632;
	 	 	 else if (in == 1323) out = -4628;
	 	 	 else if (in == 1324) out = -4625;
	 	 	 else if (in == 1325) out = -4622;
	 	 	 else if (in == 1326) out = -4619;
	 	 	 else if (in == 1327) out = -4616;
	 	 	 else if (in == 1328) out = -4613;
	 	 	 else if (in == 1329) out = -4610;
	 	 	 else if (in == 1330) out = -4607;
	 	 	 else if (in == 1331) out = -4604;
	 	 	 else if (in == 1332) out = -4601;
	 	 	 else if (in == 1333) out = -4598;
	 	 	 else if (in == 1334) out = -4595;
	 	 	 else if (in == 1335) out = -4591;
	 	 	 else if (in == 1336) out = -4588;
	 	 	 else if (in == 1337) out = -4585;
	 	 	 else if (in == 1338) out = -4582;
	 	 	 else if (in == 1339) out = -4579;
	 	 	 else if (in == 1340) out = -4576;
	 	 	 else if (in == 1341) out = -4573;
	 	 	 else if (in == 1342) out = -4570;
	 	 	 else if (in == 1343) out = -4567;
	 	 	 else if (in == 1344) out = -4564;
	 	 	 else if (in == 1345) out = -4561;
	 	 	 else if (in == 1346) out = -4558;
	 	 	 else if (in == 1347) out = -4555;
	 	 	 else if (in == 1348) out = -4552;
	 	 	 else if (in == 1349) out = -4549;
	 	 	 else if (in == 1350) out = -4546;
	 	 	 else if (in == 1351) out = -4543;
	 	 	 else if (in == 1352) out = -4540;
	 	 	 else if (in == 1353) out = -4537;
	 	 	 else if (in == 1354) out = -4534;
	 	 	 else if (in == 1355) out = -4531;
	 	 	 else if (in == 1356) out = -4528;
	 	 	 else if (in == 1357) out = -4524;
	 	 	 else if (in == 1358) out = -4521;
	 	 	 else if (in == 1359) out = -4518;
	 	 	 else if (in == 1360) out = -4515;
	 	 	 else if (in == 1361) out = -4512;
	 	 	 else if (in == 1362) out = -4509;
	 	 	 else if (in == 1363) out = -4506;
	 	 	 else if (in == 1364) out = -4503;
	 	 	 else if (in == 1365) out = -4500;
	 	 	 else if (in == 1366) out = -4497;
	 	 	 else if (in == 1367) out = -4494;
	 	 	 else if (in == 1368) out = -4491;
	 	 	 else if (in == 1369) out = -4488;
	 	 	 else if (in == 1370) out = -4485;
	 	 	 else if (in == 1371) out = -4482;
	 	 	 else if (in == 1372) out = -4479;
	 	 	 else if (in == 1373) out = -4476;
	 	 	 else if (in == 1374) out = -4473;
	 	 	 else if (in == 1375) out = -4471;
	 	 	 else if (in == 1376) out = -4468;
	 	 	 else if (in == 1377) out = -4465;
	 	 	 else if (in == 1378) out = -4462;
	 	 	 else if (in == 1379) out = -4459;
	 	 	 else if (in == 1380) out = -4456;
	 	 	 else if (in == 1381) out = -4453;
	 	 	 else if (in == 1382) out = -4450;
	 	 	 else if (in == 1383) out = -4447;
	 	 	 else if (in == 1384) out = -4444;
	 	 	 else if (in == 1385) out = -4441;
	 	 	 else if (in == 1386) out = -4438;
	 	 	 else if (in == 1387) out = -4435;
	 	 	 else if (in == 1388) out = -4432;
	 	 	 else if (in == 1389) out = -4429;
	 	 	 else if (in == 1390) out = -4426;
	 	 	 else if (in == 1391) out = -4423;
	 	 	 else if (in == 1392) out = -4420;
	 	 	 else if (in == 1393) out = -4417;
	 	 	 else if (in == 1394) out = -4414;
	 	 	 else if (in == 1395) out = -4411;
	 	 	 else if (in == 1396) out = -4408;
	 	 	 else if (in == 1397) out = -4406;
	 	 	 else if (in == 1398) out = -4403;
	 	 	 else if (in == 1399) out = -4400;
	 	 	 else if (in == 1400) out = -4397;
	 	 	 else if (in == 1401) out = -4394;
	 	 	 else if (in == 1402) out = -4391;
	 	 	 else if (in == 1403) out = -4388;
	 	 	 else if (in == 1404) out = -4385;
	 	 	 else if (in == 1405) out = -4382;
	 	 	 else if (in == 1406) out = -4379;
	 	 	 else if (in == 1407) out = -4376;
	 	 	 else if (in == 1408) out = -4373;
	 	 	 else if (in == 1409) out = -4370;
	 	 	 else if (in == 1410) out = -4368;
	 	 	 else if (in == 1411) out = -4365;
	 	 	 else if (in == 1412) out = -4362;
	 	 	 else if (in == 1413) out = -4359;
	 	 	 else if (in == 1414) out = -4356;
	 	 	 else if (in == 1415) out = -4353;
	 	 	 else if (in == 1416) out = -4350;
	 	 	 else if (in == 1417) out = -4347;
	 	 	 else if (in == 1418) out = -4344;
	 	 	 else if (in == 1419) out = -4341;
	 	 	 else if (in == 1420) out = -4339;
	 	 	 else if (in == 1421) out = -4336;
	 	 	 else if (in == 1422) out = -4333;
	 	 	 else if (in == 1423) out = -4330;
	 	 	 else if (in == 1424) out = -4327;
	 	 	 else if (in == 1425) out = -4324;
	 	 	 else if (in == 1426) out = -4321;
	 	 	 else if (in == 1427) out = -4318;
	 	 	 else if (in == 1428) out = -4316;
	 	 	 else if (in == 1429) out = -4313;
	 	 	 else if (in == 1430) out = -4310;
	 	 	 else if (in == 1431) out = -4307;
	 	 	 else if (in == 1432) out = -4304;
	 	 	 else if (in == 1433) out = -4301;
	 	 	 else if (in == 1434) out = -4298;
	 	 	 else if (in == 1435) out = -4296;
	 	 	 else if (in == 1436) out = -4293;
	 	 	 else if (in == 1437) out = -4290;
	 	 	 else if (in == 1438) out = -4287;
	 	 	 else if (in == 1439) out = -4284;
	 	 	 else if (in == 1440) out = -4281;
	 	 	 else if (in == 1441) out = -4278;
	 	 	 else if (in == 1442) out = -4276;
	 	 	 else if (in == 1443) out = -4273;
	 	 	 else if (in == 1444) out = -4270;
	 	 	 else if (in == 1445) out = -4267;
	 	 	 else if (in == 1446) out = -4264;
	 	 	 else if (in == 1447) out = -4261;
	 	 	 else if (in == 1448) out = -4259;
	 	 	 else if (in == 1449) out = -4256;
	 	 	 else if (in == 1450) out = -4253;
	 	 	 else if (in == 1451) out = -4250;
	 	 	 else if (in == 1452) out = -4247;
	 	 	 else if (in == 1453) out = -4245;
	 	 	 else if (in == 1454) out = -4242;
	 	 	 else if (in == 1455) out = -4239;
	 	 	 else if (in == 1456) out = -4236;
	 	 	 else if (in == 1457) out = -4233;
	 	 	 else if (in == 1458) out = -4230;
	 	 	 else if (in == 1459) out = -4228;
	 	 	 else if (in == 1460) out = -4225;
	 	 	 else if (in == 1461) out = -4222;
	 	 	 else if (in == 1462) out = -4219;
	 	 	 else if (in == 1463) out = -4216;
	 	 	 else if (in == 1464) out = -4214;
	 	 	 else if (in == 1465) out = -4211;
	 	 	 else if (in == 1466) out = -4208;
	 	 	 else if (in == 1467) out = -4205;
	 	 	 else if (in == 1468) out = -4202;
	 	 	 else if (in == 1469) out = -4200;
	 	 	 else if (in == 1470) out = -4197;
	 	 	 else if (in == 1471) out = -4194;
	 	 	 else if (in == 1472) out = -4191;
	 	 	 else if (in == 1473) out = -4189;
	 	 	 else if (in == 1474) out = -4186;
	 	 	 else if (in == 1475) out = -4183;
	 	 	 else if (in == 1476) out = -4180;
	 	 	 else if (in == 1477) out = -4177;
	 	 	 else if (in == 1478) out = -4175;
	 	 	 else if (in == 1479) out = -4172;
	 	 	 else if (in == 1480) out = -4169;
	 	 	 else if (in == 1481) out = -4166;
	 	 	 else if (in == 1482) out = -4164;
	 	 	 else if (in == 1483) out = -4161;
	 	 	 else if (in == 1484) out = -4158;
	 	 	 else if (in == 1485) out = -4155;
	 	 	 else if (in == 1486) out = -4153;
	 	 	 else if (in == 1487) out = -4150;
	 	 	 else if (in == 1488) out = -4147;
	 	 	 else if (in == 1489) out = -4144;
	 	 	 else if (in == 1490) out = -4142;
	 	 	 else if (in == 1491) out = -4139;
	 	 	 else if (in == 1492) out = -4136;
	 	 	 else if (in == 1493) out = -4133;
	 	 	 else if (in == 1494) out = -4131;
	 	 	 else if (in == 1495) out = -4128;
	 	 	 else if (in == 1496) out = -4125;
	 	 	 else if (in == 1497) out = -4122;
	 	 	 else if (in == 1498) out = -4120;
	 	 	 else if (in == 1499) out = -4117;
	 	 	 else if (in == 1500) out = -4114;
	 	 	 else if (in == 1501) out = -4111;
	 	 	 else if (in == 1502) out = -4109;
	 	 	 else if (in == 1503) out = -4106;
	 	 	 else if (in == 1504) out = -4103;
	 	 	 else if (in == 1505) out = -4100;
	 	 	 else if (in == 1506) out = -4098;
	 	 	 else if (in == 1507) out = -4095;
	 	 	 else if (in == 1508) out = -4092;
	 	 	 else if (in == 1509) out = -4090;
	 	 	 else if (in == 1510) out = -4087;
	 	 	 else if (in == 1511) out = -4084;
	 	 	 else if (in == 1512) out = -4081;
	 	 	 else if (in == 1513) out = -4079;
	 	 	 else if (in == 1514) out = -4076;
	 	 	 else if (in == 1515) out = -4073;
	 	 	 else if (in == 1516) out = -4071;
	 	 	 else if (in == 1517) out = -4068;
	 	 	 else if (in == 1518) out = -4065;
	 	 	 else if (in == 1519) out = -4063;
	 	 	 else if (in == 1520) out = -4060;
	 	 	 else if (in == 1521) out = -4057;
	 	 	 else if (in == 1522) out = -4054;
	 	 	 else if (in == 1523) out = -4052;
	 	 	 else if (in == 1524) out = -4049;
	 	 	 else if (in == 1525) out = -4046;
	 	 	 else if (in == 1526) out = -4044;
	 	 	 else if (in == 1527) out = -4041;
	 	 	 else if (in == 1528) out = -4038;
	 	 	 else if (in == 1529) out = -4036;
	 	 	 else if (in == 1530) out = -4033;
	 	 	 else if (in == 1531) out = -4030;
	 	 	 else if (in == 1532) out = -4028;
	 	 	 else if (in == 1533) out = -4025;
	 	 	 else if (in == 1534) out = -4022;
	 	 	 else if (in == 1535) out = -4020;
	 	 	 else if (in == 1536) out = -4017;
	 	 	 else if (in == 1537) out = -4014;
	 	 	 else if (in == 1538) out = -4012;
	 	 	 else if (in == 1539) out = -4009;
	 	 	 else if (in == 1540) out = -4006;
	 	 	 else if (in == 1541) out = -4004;
	 	 	 else if (in == 1542) out = -4001;
	 	 	 else if (in == 1543) out = -3998;
	 	 	 else if (in == 1544) out = -3996;
	 	 	 else if (in == 1545) out = -3993;
	 	 	 else if (in == 1546) out = -3990;
	 	 	 else if (in == 1547) out = -3988;
	 	 	 else if (in == 1548) out = -3985;
	 	 	 else if (in == 1549) out = -3982;
	 	 	 else if (in == 1550) out = -3980;
	 	 	 else if (in == 1551) out = -3977;
	 	 	 else if (in == 1552) out = -3975;
	 	 	 else if (in == 1553) out = -3972;
	 	 	 else if (in == 1554) out = -3969;
	 	 	 else if (in == 1555) out = -3967;
	 	 	 else if (in == 1556) out = -3964;
	 	 	 else if (in == 1557) out = -3961;
	 	 	 else if (in == 1558) out = -3959;
	 	 	 else if (in == 1559) out = -3956;
	 	 	 else if (in == 1560) out = -3953;
	 	 	 else if (in == 1561) out = -3951;
	 	 	 else if (in == 1562) out = -3948;
	 	 	 else if (in == 1563) out = -3946;
	 	 	 else if (in == 1564) out = -3943;
	 	 	 else if (in == 1565) out = -3940;
	 	 	 else if (in == 1566) out = -3938;
	 	 	 else if (in == 1567) out = -3935;
	 	 	 else if (in == 1568) out = -3933;
	 	 	 else if (in == 1569) out = -3930;
	 	 	 else if (in == 1570) out = -3927;
	 	 	 else if (in == 1571) out = -3925;
	 	 	 else if (in == 1572) out = -3922;
	 	 	 else if (in == 1573) out = -3919;
	 	 	 else if (in == 1574) out = -3917;
	 	 	 else if (in == 1575) out = -3914;
	 	 	 else if (in == 1576) out = -3912;
	 	 	 else if (in == 1577) out = -3909;
	 	 	 else if (in == 1578) out = -3906;
	 	 	 else if (in == 1579) out = -3904;
	 	 	 else if (in == 1580) out = -3901;
	 	 	 else if (in == 1581) out = -3899;
	 	 	 else if (in == 1582) out = -3896;
	 	 	 else if (in == 1583) out = -3894;
	 	 	 else if (in == 1584) out = -3891;
	 	 	 else if (in == 1585) out = -3888;
	 	 	 else if (in == 1586) out = -3886;
	 	 	 else if (in == 1587) out = -3883;
	 	 	 else if (in == 1588) out = -3881;
	 	 	 else if (in == 1589) out = -3878;
	 	 	 else if (in == 1590) out = -3875;
	 	 	 else if (in == 1591) out = -3873;
	 	 	 else if (in == 1592) out = -3870;
	 	 	 else if (in == 1593) out = -3868;
	 	 	 else if (in == 1594) out = -3865;
	 	 	 else if (in == 1595) out = -3863;
	 	 	 else if (in == 1596) out = -3860;
	 	 	 else if (in == 1597) out = -3857;
	 	 	 else if (in == 1598) out = -3855;
	 	 	 else if (in == 1599) out = -3852;
	 	 	 else if (in == 1600) out = -3850;
	 	 	 else if (in == 1601) out = -3847;
	 	 	 else if (in == 1602) out = -3845;
	 	 	 else if (in == 1603) out = -3842;
	 	 	 else if (in == 1604) out = -3840;
	 	 	 else if (in == 1605) out = -3837;
	 	 	 else if (in == 1606) out = -3834;
	 	 	 else if (in == 1607) out = -3832;
	 	 	 else if (in == 1608) out = -3829;
	 	 	 else if (in == 1609) out = -3827;
	 	 	 else if (in == 1610) out = -3824;
	 	 	 else if (in == 1611) out = -3822;
	 	 	 else if (in == 1612) out = -3819;
	 	 	 else if (in == 1613) out = -3817;
	 	 	 else if (in == 1614) out = -3814;
	 	 	 else if (in == 1615) out = -3812;
	 	 	 else if (in == 1616) out = -3809;
	 	 	 else if (in == 1617) out = -3806;
	 	 	 else if (in == 1618) out = -3804;
	 	 	 else if (in == 1619) out = -3801;
	 	 	 else if (in == 1620) out = -3799;
	 	 	 else if (in == 1621) out = -3796;
	 	 	 else if (in == 1622) out = -3794;
	 	 	 else if (in == 1623) out = -3791;
	 	 	 else if (in == 1624) out = -3789;
	 	 	 else if (in == 1625) out = -3786;
	 	 	 else if (in == 1626) out = -3784;
	 	 	 else if (in == 1627) out = -3781;
	 	 	 else if (in == 1628) out = -3779;
	 	 	 else if (in == 1629) out = -3776;
	 	 	 else if (in == 1630) out = -3774;
	 	 	 else if (in == 1631) out = -3771;
	 	 	 else if (in == 1632) out = -3769;
	 	 	 else if (in == 1633) out = -3766;
	 	 	 else if (in == 1634) out = -3764;
	 	 	 else if (in == 1635) out = -3761;
	 	 	 else if (in == 1636) out = -3759;
	 	 	 else if (in == 1637) out = -3756;
	 	 	 else if (in == 1638) out = -3754;
	 	 	 else if (in == 1639) out = -3751;
	 	 	 else if (in == 1640) out = -3749;
	 	 	 else if (in == 1641) out = -3746;
	 	 	 else if (in == 1642) out = -3744;
	 	 	 else if (in == 1643) out = -3741;
	 	 	 else if (in == 1644) out = -3739;
	 	 	 else if (in == 1645) out = -3736;
	 	 	 else if (in == 1646) out = -3734;
	 	 	 else if (in == 1647) out = -3731;
	 	 	 else if (in == 1648) out = -3729;
	 	 	 else if (in == 1649) out = -3726;
	 	 	 else if (in == 1650) out = -3724;
	 	 	 else if (in == 1651) out = -3721;
	 	 	 else if (in == 1652) out = -3719;
	 	 	 else if (in == 1653) out = -3716;
	 	 	 else if (in == 1654) out = -3714;
	 	 	 else if (in == 1655) out = -3711;
	 	 	 else if (in == 1656) out = -3709;
	 	 	 else if (in == 1657) out = -3706;
	 	 	 else if (in == 1658) out = -3704;
	 	 	 else if (in == 1659) out = -3701;
	 	 	 else if (in == 1660) out = -3699;
	 	 	 else if (in == 1661) out = -3697;
	 	 	 else if (in == 1662) out = -3694;
	 	 	 else if (in == 1663) out = -3692;
	 	 	 else if (in == 1664) out = -3689;
	 	 	 else if (in == 1665) out = -3687;
	 	 	 else if (in == 1666) out = -3684;
	 	 	 else if (in == 1667) out = -3682;
	 	 	 else if (in == 1668) out = -3679;
	 	 	 else if (in == 1669) out = -3677;
	 	 	 else if (in == 1670) out = -3674;
	 	 	 else if (in == 1671) out = -3672;
	 	 	 else if (in == 1672) out = -3669;
	 	 	 else if (in == 1673) out = -3667;
	 	 	 else if (in == 1674) out = -3665;
	 	 	 else if (in == 1675) out = -3662;
	 	 	 else if (in == 1676) out = -3660;
	 	 	 else if (in == 1677) out = -3657;
	 	 	 else if (in == 1678) out = -3655;
	 	 	 else if (in == 1679) out = -3652;
	 	 	 else if (in == 1680) out = -3650;
	 	 	 else if (in == 1681) out = -3647;
	 	 	 else if (in == 1682) out = -3645;
	 	 	 else if (in == 1683) out = -3643;
	 	 	 else if (in == 1684) out = -3640;
	 	 	 else if (in == 1685) out = -3638;
	 	 	 else if (in == 1686) out = -3635;
	 	 	 else if (in == 1687) out = -3633;
	 	 	 else if (in == 1688) out = -3630;
	 	 	 else if (in == 1689) out = -3628;
	 	 	 else if (in == 1690) out = -3626;
	 	 	 else if (in == 1691) out = -3623;
	 	 	 else if (in == 1692) out = -3621;
	 	 	 else if (in == 1693) out = -3618;
	 	 	 else if (in == 1694) out = -3616;
	 	 	 else if (in == 1695) out = -3614;
	 	 	 else if (in == 1696) out = -3611;
	 	 	 else if (in == 1697) out = -3609;
	 	 	 else if (in == 1698) out = -3606;
	 	 	 else if (in == 1699) out = -3604;
	 	 	 else if (in == 1700) out = -3601;
	 	 	 else if (in == 1701) out = -3599;
	 	 	 else if (in == 1702) out = -3597;
	 	 	 else if (in == 1703) out = -3594;
	 	 	 else if (in == 1704) out = -3592;
	 	 	 else if (in == 1705) out = -3589;
	 	 	 else if (in == 1706) out = -3587;
	 	 	 else if (in == 1707) out = -3585;
	 	 	 else if (in == 1708) out = -3582;
	 	 	 else if (in == 1709) out = -3580;
	 	 	 else if (in == 1710) out = -3577;
	 	 	 else if (in == 1711) out = -3575;
	 	 	 else if (in == 1712) out = -3573;
	 	 	 else if (in == 1713) out = -3570;
	 	 	 else if (in == 1714) out = -3568;
	 	 	 else if (in == 1715) out = -3565;
	 	 	 else if (in == 1716) out = -3563;
	 	 	 else if (in == 1717) out = -3561;
	 	 	 else if (in == 1718) out = -3558;
	 	 	 else if (in == 1719) out = -3556;
	 	 	 else if (in == 1720) out = -3554;
	 	 	 else if (in == 1721) out = -3551;
	 	 	 else if (in == 1722) out = -3549;
	 	 	 else if (in == 1723) out = -3546;
	 	 	 else if (in == 1724) out = -3544;
	 	 	 else if (in == 1725) out = -3542;
	 	 	 else if (in == 1726) out = -3539;
	 	 	 else if (in == 1727) out = -3537;
	 	 	 else if (in == 1728) out = -3535;
	 	 	 else if (in == 1729) out = -3532;
	 	 	 else if (in == 1730) out = -3530;
	 	 	 else if (in == 1731) out = -3527;
	 	 	 else if (in == 1732) out = -3525;
	 	 	 else if (in == 1733) out = -3523;
	 	 	 else if (in == 1734) out = -3520;
	 	 	 else if (in == 1735) out = -3518;
	 	 	 else if (in == 1736) out = -3516;
	 	 	 else if (in == 1737) out = -3513;
	 	 	 else if (in == 1738) out = -3511;
	 	 	 else if (in == 1739) out = -3509;
	 	 	 else if (in == 1740) out = -3506;
	 	 	 else if (in == 1741) out = -3504;
	 	 	 else if (in == 1742) out = -3501;
	 	 	 else if (in == 1743) out = -3499;
	 	 	 else if (in == 1744) out = -3497;
	 	 	 else if (in == 1745) out = -3494;
	 	 	 else if (in == 1746) out = -3492;
	 	 	 else if (in == 1747) out = -3490;
	 	 	 else if (in == 1748) out = -3487;
	 	 	 else if (in == 1749) out = -3485;
	 	 	 else if (in == 1750) out = -3483;
	 	 	 else if (in == 1751) out = -3480;
	 	 	 else if (in == 1752) out = -3478;
	 	 	 else if (in == 1753) out = -3476;
	 	 	 else if (in == 1754) out = -3473;
	 	 	 else if (in == 1755) out = -3471;
	 	 	 else if (in == 1756) out = -3469;
	 	 	 else if (in == 1757) out = -3466;
	 	 	 else if (in == 1758) out = -3464;
	 	 	 else if (in == 1759) out = -3462;
	 	 	 else if (in == 1760) out = -3459;
	 	 	 else if (in == 1761) out = -3457;
	 	 	 else if (in == 1762) out = -3455;
	 	 	 else if (in == 1763) out = -3452;
	 	 	 else if (in == 1764) out = -3450;
	 	 	 else if (in == 1765) out = -3448;
	 	 	 else if (in == 1766) out = -3445;
	 	 	 else if (in == 1767) out = -3443;
	 	 	 else if (in == 1768) out = -3441;
	 	 	 else if (in == 1769) out = -3438;
	 	 	 else if (in == 1770) out = -3436;
	 	 	 else if (in == 1771) out = -3434;
	 	 	 else if (in == 1772) out = -3432;
	 	 	 else if (in == 1773) out = -3429;
	 	 	 else if (in == 1774) out = -3427;
	 	 	 else if (in == 1775) out = -3425;
	 	 	 else if (in == 1776) out = -3422;
	 	 	 else if (in == 1777) out = -3420;
	 	 	 else if (in == 1778) out = -3418;
	 	 	 else if (in == 1779) out = -3415;
	 	 	 else if (in == 1780) out = -3413;
	 	 	 else if (in == 1781) out = -3411;
	 	 	 else if (in == 1782) out = -3408;
	 	 	 else if (in == 1783) out = -3406;
	 	 	 else if (in == 1784) out = -3404;
	 	 	 else if (in == 1785) out = -3402;
	 	 	 else if (in == 1786) out = -3399;
	 	 	 else if (in == 1787) out = -3397;
	 	 	 else if (in == 1788) out = -3395;
	 	 	 else if (in == 1789) out = -3392;
	 	 	 else if (in == 1790) out = -3390;
	 	 	 else if (in == 1791) out = -3388;
	 	 	 else if (in == 1792) out = -3386;
	 	 	 else if (in == 1793) out = -3383;
	 	 	 else if (in == 1794) out = -3381;
	 	 	 else if (in == 1795) out = -3379;
	 	 	 else if (in == 1796) out = -3376;
	 	 	 else if (in == 1797) out = -3374;
	 	 	 else if (in == 1798) out = -3372;
	 	 	 else if (in == 1799) out = -3370;
	 	 	 else if (in == 1800) out = -3367;
	 	 	 else if (in == 1801) out = -3365;
	 	 	 else if (in == 1802) out = -3363;
	 	 	 else if (in == 1803) out = -3361;
	 	 	 else if (in == 1804) out = -3358;
	 	 	 else if (in == 1805) out = -3356;
	 	 	 else if (in == 1806) out = -3354;
	 	 	 else if (in == 1807) out = -3351;
	 	 	 else if (in == 1808) out = -3349;
	 	 	 else if (in == 1809) out = -3347;
	 	 	 else if (in == 1810) out = -3345;
	 	 	 else if (in == 1811) out = -3342;
	 	 	 else if (in == 1812) out = -3340;
	 	 	 else if (in == 1813) out = -3338;
	 	 	 else if (in == 1814) out = -3336;
	 	 	 else if (in == 1815) out = -3333;
	 	 	 else if (in == 1816) out = -3331;
	 	 	 else if (in == 1817) out = -3329;
	 	 	 else if (in == 1818) out = -3327;
	 	 	 else if (in == 1819) out = -3324;
	 	 	 else if (in == 1820) out = -3322;
	 	 	 else if (in == 1821) out = -3320;
	 	 	 else if (in == 1822) out = -3318;
	 	 	 else if (in == 1823) out = -3315;
	 	 	 else if (in == 1824) out = -3313;
	 	 	 else if (in == 1825) out = -3311;
	 	 	 else if (in == 1826) out = -3309;
	 	 	 else if (in == 1827) out = -3306;
	 	 	 else if (in == 1828) out = -3304;
	 	 	 else if (in == 1829) out = -3302;
	 	 	 else if (in == 1830) out = -3300;
	 	 	 else if (in == 1831) out = -3297;
	 	 	 else if (in == 1832) out = -3295;
	 	 	 else if (in == 1833) out = -3293;
	 	 	 else if (in == 1834) out = -3291;
	 	 	 else if (in == 1835) out = -3288;
	 	 	 else if (in == 1836) out = -3286;
	 	 	 else if (in == 1837) out = -3284;
	 	 	 else if (in == 1838) out = -3282;
	 	 	 else if (in == 1839) out = -3280;
	 	 	 else if (in == 1840) out = -3277;
	 	 	 else if (in == 1841) out = -3275;
	 	 	 else if (in == 1842) out = -3273;
	 	 	 else if (in == 1843) out = -3271;
	 	 	 else if (in == 1844) out = -3268;
	 	 	 else if (in == 1845) out = -3266;
	 	 	 else if (in == 1846) out = -3264;
	 	 	 else if (in == 1847) out = -3262;
	 	 	 else if (in == 1848) out = -3260;
	 	 	 else if (in == 1849) out = -3257;
	 	 	 else if (in == 1850) out = -3255;
	 	 	 else if (in == 1851) out = -3253;
	 	 	 else if (in == 1852) out = -3251;
	 	 	 else if (in == 1853) out = -3248;
	 	 	 else if (in == 1854) out = -3246;
	 	 	 else if (in == 1855) out = -3244;
	 	 	 else if (in == 1856) out = -3242;
	 	 	 else if (in == 1857) out = -3240;
	 	 	 else if (in == 1858) out = -3237;
	 	 	 else if (in == 1859) out = -3235;
	 	 	 else if (in == 1860) out = -3233;
	 	 	 else if (in == 1861) out = -3231;
	 	 	 else if (in == 1862) out = -3229;
	 	 	 else if (in == 1863) out = -3226;
	 	 	 else if (in == 1864) out = -3224;
	 	 	 else if (in == 1865) out = -3222;
	 	 	 else if (in == 1866) out = -3220;
	 	 	 else if (in == 1867) out = -3218;
	 	 	 else if (in == 1868) out = -3215;
	 	 	 else if (in == 1869) out = -3213;
	 	 	 else if (in == 1870) out = -3211;
	 	 	 else if (in == 1871) out = -3209;
	 	 	 else if (in == 1872) out = -3207;
	 	 	 else if (in == 1873) out = -3204;
	 	 	 else if (in == 1874) out = -3202;
	 	 	 else if (in == 1875) out = -3200;
	 	 	 else if (in == 1876) out = -3198;
	 	 	 else if (in == 1877) out = -3196;
	 	 	 else if (in == 1878) out = -3194;
	 	 	 else if (in == 1879) out = -3191;
	 	 	 else if (in == 1880) out = -3189;
	 	 	 else if (in == 1881) out = -3187;
	 	 	 else if (in == 1882) out = -3185;
	 	 	 else if (in == 1883) out = -3183;
	 	 	 else if (in == 1884) out = -3181;
	 	 	 else if (in == 1885) out = -3178;
	 	 	 else if (in == 1886) out = -3176;
	 	 	 else if (in == 1887) out = -3174;
	 	 	 else if (in == 1888) out = -3172;
	 	 	 else if (in == 1889) out = -3170;
	 	 	 else if (in == 1890) out = -3167;
	 	 	 else if (in == 1891) out = -3165;
	 	 	 else if (in == 1892) out = -3163;
	 	 	 else if (in == 1893) out = -3161;
	 	 	 else if (in == 1894) out = -3159;
	 	 	 else if (in == 1895) out = -3157;
	 	 	 else if (in == 1896) out = -3155;
	 	 	 else if (in == 1897) out = -3152;
	 	 	 else if (in == 1898) out = -3150;
	 	 	 else if (in == 1899) out = -3148;
	 	 	 else if (in == 1900) out = -3146;
	 	 	 else if (in == 1901) out = -3144;
	 	 	 else if (in == 1902) out = -3142;
	 	 	 else if (in == 1903) out = -3139;
	 	 	 else if (in == 1904) out = -3137;
	 	 	 else if (in == 1905) out = -3135;
	 	 	 else if (in == 1906) out = -3133;
	 	 	 else if (in == 1907) out = -3131;
	 	 	 else if (in == 1908) out = -3129;
	 	 	 else if (in == 1909) out = -3127;
	 	 	 else if (in == 1910) out = -3124;
	 	 	 else if (in == 1911) out = -3122;
	 	 	 else if (in == 1912) out = -3120;
	 	 	 else if (in == 1913) out = -3118;
	 	 	 else if (in == 1914) out = -3116;
	 	 	 else if (in == 1915) out = -3114;
	 	 	 else if (in == 1916) out = -3112;
	 	 	 else if (in == 1917) out = -3109;
	 	 	 else if (in == 1918) out = -3107;
	 	 	 else if (in == 1919) out = -3105;
	 	 	 else if (in == 1920) out = -3103;
	 	 	 else if (in == 1921) out = -3101;
	 	 	 else if (in == 1922) out = -3099;
	 	 	 else if (in == 1923) out = -3097;
	 	 	 else if (in == 1924) out = -3094;
	 	 	 else if (in == 1925) out = -3092;
	 	 	 else if (in == 1926) out = -3090;
	 	 	 else if (in == 1927) out = -3088;
	 	 	 else if (in == 1928) out = -3086;
	 	 	 else if (in == 1929) out = -3084;
	 	 	 else if (in == 1930) out = -3082;
	 	 	 else if (in == 1931) out = -3080;
	 	 	 else if (in == 1932) out = -3077;
	 	 	 else if (in == 1933) out = -3075;
	 	 	 else if (in == 1934) out = -3073;
	 	 	 else if (in == 1935) out = -3071;
	 	 	 else if (in == 1936) out = -3069;
	 	 	 else if (in == 1937) out = -3067;
	 	 	 else if (in == 1938) out = -3065;
	 	 	 else if (in == 1939) out = -3063;
	 	 	 else if (in == 1940) out = -3061;
	 	 	 else if (in == 1941) out = -3058;
	 	 	 else if (in == 1942) out = -3056;
	 	 	 else if (in == 1943) out = -3054;
	 	 	 else if (in == 1944) out = -3052;
	 	 	 else if (in == 1945) out = -3050;
	 	 	 else if (in == 1946) out = -3048;
	 	 	 else if (in == 1947) out = -3046;
	 	 	 else if (in == 1948) out = -3044;
	 	 	 else if (in == 1949) out = -3042;
	 	 	 else if (in == 1950) out = -3039;
	 	 	 else if (in == 1951) out = -3037;
	 	 	 else if (in == 1952) out = -3035;
	 	 	 else if (in == 1953) out = -3033;
	 	 	 else if (in == 1954) out = -3031;
	 	 	 else if (in == 1955) out = -3029;
	 	 	 else if (in == 1956) out = -3027;
	 	 	 else if (in == 1957) out = -3025;
	 	 	 else if (in == 1958) out = -3023;
	 	 	 else if (in == 1959) out = -3021;
	 	 	 else if (in == 1960) out = -3019;
	 	 	 else if (in == 1961) out = -3016;
	 	 	 else if (in == 1962) out = -3014;
	 	 	 else if (in == 1963) out = -3012;
	 	 	 else if (in == 1964) out = -3010;
	 	 	 else if (in == 1965) out = -3008;
	 	 	 else if (in == 1966) out = -3006;
	 	 	 else if (in == 1967) out = -3004;
	 	 	 else if (in == 1968) out = -3002;
	 	 	 else if (in == 1969) out = -3000;
	 	 	 else if (in == 1970) out = -2998;
	 	 	 else if (in == 1971) out = -2996;
	 	 	 else if (in == 1972) out = -2994;
	 	 	 else if (in == 1973) out = -2991;
	 	 	 else if (in == 1974) out = -2989;
	 	 	 else if (in == 1975) out = -2987;
	 	 	 else if (in == 1976) out = -2985;
	 	 	 else if (in == 1977) out = -2983;
	 	 	 else if (in == 1978) out = -2981;
	 	 	 else if (in == 1979) out = -2979;
	 	 	 else if (in == 1980) out = -2977;
	 	 	 else if (in == 1981) out = -2975;
	 	 	 else if (in == 1982) out = -2973;
	 	 	 else if (in == 1983) out = -2971;
	 	 	 else if (in == 1984) out = -2969;
	 	 	 else if (in == 1985) out = -2967;
	 	 	 else if (in == 1986) out = -2965;
	 	 	 else if (in == 1987) out = -2962;
	 	 	 else if (in == 1988) out = -2960;
	 	 	 else if (in == 1989) out = -2958;
	 	 	 else if (in == 1990) out = -2956;
	 	 	 else if (in == 1991) out = -2954;
	 	 	 else if (in == 1992) out = -2952;
	 	 	 else if (in == 1993) out = -2950;
	 	 	 else if (in == 1994) out = -2948;
	 	 	 else if (in == 1995) out = -2946;
	 	 	 else if (in == 1996) out = -2944;
	 	 	 else if (in == 1997) out = -2942;
	 	 	 else if (in == 1998) out = -2940;
	 	 	 else if (in == 1999) out = -2938;
	 	 	 else if (in == 2000) out = -2936;
	 	 	 else if (in == 2001) out = -2934;
	 	 	 else if (in == 2002) out = -2932;
	 	 	 else if (in == 2003) out = -2930;
	 	 	 else if (in == 2004) out = -2928;
	 	 	 else if (in == 2005) out = -2926;
	 	 	 else if (in == 2006) out = -2924;
	 	 	 else if (in == 2007) out = -2921;
	 	 	 else if (in == 2008) out = -2919;
	 	 	 else if (in == 2009) out = -2917;
	 	 	 else if (in == 2010) out = -2915;
	 	 	 else if (in == 2011) out = -2913;
	 	 	 else if (in == 2012) out = -2911;
	 	 	 else if (in == 2013) out = -2909;
	 	 	 else if (in == 2014) out = -2907;
	 	 	 else if (in == 2015) out = -2905;
	 	 	 else if (in == 2016) out = -2903;
	 	 	 else if (in == 2017) out = -2901;
	 	 	 else if (in == 2018) out = -2899;
	 	 	 else if (in == 2019) out = -2897;
	 	 	 else if (in == 2020) out = -2895;
	 	 	 else if (in == 2021) out = -2893;
	 	 	 else if (in == 2022) out = -2891;
	 	 	 else if (in == 2023) out = -2889;
	 	 	 else if (in == 2024) out = -2887;
	 	 	 else if (in == 2025) out = -2885;
	 	 	 else if (in == 2026) out = -2883;
	 	 	 else if (in == 2027) out = -2881;
	 	 	 else if (in == 2028) out = -2879;
	 	 	 else if (in == 2029) out = -2877;
	 	 	 else if (in == 2030) out = -2875;
	 	 	 else if (in == 2031) out = -2873;
	 	 	 else if (in == 2032) out = -2871;
	 	 	 else if (in == 2033) out = -2869;
	 	 	 else if (in == 2034) out = -2867;
	 	 	 else if (in == 2035) out = -2865;
	 	 	 else if (in == 2036) out = -2863;
	 	 	 else if (in == 2037) out = -2861;
	 	 	 else if (in == 2038) out = -2859;
	 	 	 else if (in == 2039) out = -2857;
	 	 	 else if (in == 2040) out = -2855;
	 	 	 else if (in == 2041) out = -2853;
	 	 	 else if (in == 2042) out = -2851;
	 	 	 else if (in == 2043) out = -2849;
	 	 	 else if (in == 2044) out = -2847;
	 	 	 else if (in == 2045) out = -2845;
	 	 	 else if (in == 2046) out = -2843;
	 	 	 else if (in == 2047) out = -2841;
	 	 	 else if (in == 2048) out = -2839;
	 	 	 else if (in == 2049) out = -2837;
	 	 	 else if (in == 2050) out = -2835;
	 	 	 else if (in == 2051) out = -2833;
	 	 	 else if (in == 2052) out = -2831;
	 	 	 else if (in == 2053) out = -2829;
	 	 	 else if (in == 2054) out = -2827;
	 	 	 else if (in == 2055) out = -2825;
	 	 	 else if (in == 2056) out = -2823;
	 	 	 else if (in == 2057) out = -2821;
	 	 	 else if (in == 2058) out = -2819;
	 	 	 else if (in == 2059) out = -2817;
	 	 	 else if (in == 2060) out = -2815;
	 	 	 else if (in == 2061) out = -2813;
	 	 	 else if (in == 2062) out = -2811;
	 	 	 else if (in == 2063) out = -2809;
	 	 	 else if (in == 2064) out = -2807;
	 	 	 else if (in == 2065) out = -2805;
	 	 	 else if (in == 2066) out = -2803;
	 	 	 else if (in == 2067) out = -2801;
	 	 	 else if (in == 2068) out = -2799;
	 	 	 else if (in == 2069) out = -2797;
	 	 	 else if (in == 2070) out = -2795;
	 	 	 else if (in == 2071) out = -2793;
	 	 	 else if (in == 2072) out = -2791;
	 	 	 else if (in == 2073) out = -2789;
	 	 	 else if (in == 2074) out = -2787;
	 	 	 else if (in == 2075) out = -2785;
	 	 	 else if (in == 2076) out = -2783;
	 	 	 else if (in == 2077) out = -2781;
	 	 	 else if (in == 2078) out = -2779;
	 	 	 else if (in == 2079) out = -2777;
	 	 	 else if (in == 2080) out = -2775;
	 	 	 else if (in == 2081) out = -2773;
	 	 	 else if (in == 2082) out = -2771;
	 	 	 else if (in == 2083) out = -2769;
	 	 	 else if (in == 2084) out = -2767;
	 	 	 else if (in == 2085) out = -2765;
	 	 	 else if (in == 2086) out = -2763;
	 	 	 else if (in == 2087) out = -2761;
	 	 	 else if (in == 2088) out = -2759;
	 	 	 else if (in == 2089) out = -2757;
	 	 	 else if (in == 2090) out = -2755;
	 	 	 else if (in == 2091) out = -2754;
	 	 	 else if (in == 2092) out = -2752;
	 	 	 else if (in == 2093) out = -2750;
	 	 	 else if (in == 2094) out = -2748;
	 	 	 else if (in == 2095) out = -2746;
	 	 	 else if (in == 2096) out = -2744;
	 	 	 else if (in == 2097) out = -2742;
	 	 	 else if (in == 2098) out = -2740;
	 	 	 else if (in == 2099) out = -2738;
	 	 	 else if (in == 2100) out = -2736;
	 	 	 else if (in == 2101) out = -2734;
	 	 	 else if (in == 2102) out = -2732;
	 	 	 else if (in == 2103) out = -2730;
	 	 	 else if (in == 2104) out = -2728;
	 	 	 else if (in == 2105) out = -2726;
	 	 	 else if (in == 2106) out = -2724;
	 	 	 else if (in == 2107) out = -2722;
	 	 	 else if (in == 2108) out = -2720;
	 	 	 else if (in == 2109) out = -2718;
	 	 	 else if (in == 2110) out = -2716;
	 	 	 else if (in == 2111) out = -2715;
	 	 	 else if (in == 2112) out = -2713;
	 	 	 else if (in == 2113) out = -2711;
	 	 	 else if (in == 2114) out = -2709;
	 	 	 else if (in == 2115) out = -2707;
	 	 	 else if (in == 2116) out = -2705;
	 	 	 else if (in == 2117) out = -2703;
	 	 	 else if (in == 2118) out = -2701;
	 	 	 else if (in == 2119) out = -2699;
	 	 	 else if (in == 2120) out = -2697;
	 	 	 else if (in == 2121) out = -2695;
	 	 	 else if (in == 2122) out = -2693;
	 	 	 else if (in == 2123) out = -2691;
	 	 	 else if (in == 2124) out = -2689;
	 	 	 else if (in == 2125) out = -2687;
	 	 	 else if (in == 2126) out = -2686;
	 	 	 else if (in == 2127) out = -2684;
	 	 	 else if (in == 2128) out = -2682;
	 	 	 else if (in == 2129) out = -2680;
	 	 	 else if (in == 2130) out = -2678;
	 	 	 else if (in == 2131) out = -2676;
	 	 	 else if (in == 2132) out = -2674;
	 	 	 else if (in == 2133) out = -2672;
	 	 	 else if (in == 2134) out = -2670;
	 	 	 else if (in == 2135) out = -2668;
	 	 	 else if (in == 2136) out = -2666;
	 	 	 else if (in == 2137) out = -2664;
	 	 	 else if (in == 2138) out = -2662;
	 	 	 else if (in == 2139) out = -2661;
	 	 	 else if (in == 2140) out = -2659;
	 	 	 else if (in == 2141) out = -2657;
	 	 	 else if (in == 2142) out = -2655;
	 	 	 else if (in == 2143) out = -2653;
	 	 	 else if (in == 2144) out = -2651;
	 	 	 else if (in == 2145) out = -2649;
	 	 	 else if (in == 2146) out = -2647;
	 	 	 else if (in == 2147) out = -2645;
	 	 	 else if (in == 2148) out = -2643;
	 	 	 else if (in == 2149) out = -2641;
	 	 	 else if (in == 2150) out = -2640;
	 	 	 else if (in == 2151) out = -2638;
	 	 	 else if (in == 2152) out = -2636;
	 	 	 else if (in == 2153) out = -2634;
	 	 	 else if (in == 2154) out = -2632;
	 	 	 else if (in == 2155) out = -2630;
	 	 	 else if (in == 2156) out = -2628;
	 	 	 else if (in == 2157) out = -2626;
	 	 	 else if (in == 2158) out = -2624;
	 	 	 else if (in == 2159) out = -2622;
	 	 	 else if (in == 2160) out = -2621;
	 	 	 else if (in == 2161) out = -2619;
	 	 	 else if (in == 2162) out = -2617;
	 	 	 else if (in == 2163) out = -2615;
	 	 	 else if (in == 2164) out = -2613;
	 	 	 else if (in == 2165) out = -2611;
	 	 	 else if (in == 2166) out = -2609;
	 	 	 else if (in == 2167) out = -2607;
	 	 	 else if (in == 2168) out = -2605;
	 	 	 else if (in == 2169) out = -2604;
	 	 	 else if (in == 2170) out = -2602;
	 	 	 else if (in == 2171) out = -2600;
	 	 	 else if (in == 2172) out = -2598;
	 	 	 else if (in == 2173) out = -2596;
	 	 	 else if (in == 2174) out = -2594;
	 	 	 else if (in == 2175) out = -2592;
	 	 	 else if (in == 2176) out = -2590;
	 	 	 else if (in == 2177) out = -2588;
	 	 	 else if (in == 2178) out = -2587;
	 	 	 else if (in == 2179) out = -2585;
	 	 	 else if (in == 2180) out = -2583;
	 	 	 else if (in == 2181) out = -2581;
	 	 	 else if (in == 2182) out = -2579;
	 	 	 else if (in == 2183) out = -2577;
	 	 	 else if (in == 2184) out = -2575;
	 	 	 else if (in == 2185) out = -2573;
	 	 	 else if (in == 2186) out = -2572;
	 	 	 else if (in == 2187) out = -2570;
	 	 	 else if (in == 2188) out = -2568;
	 	 	 else if (in == 2189) out = -2566;
	 	 	 else if (in == 2190) out = -2564;
	 	 	 else if (in == 2191) out = -2562;
	 	 	 else if (in == 2192) out = -2560;
	 	 	 else if (in == 2193) out = -2558;
	 	 	 else if (in == 2194) out = -2557;
	 	 	 else if (in == 2195) out = -2555;
	 	 	 else if (in == 2196) out = -2553;
	 	 	 else if (in == 2197) out = -2551;
	 	 	 else if (in == 2198) out = -2549;
	 	 	 else if (in == 2199) out = -2547;
	 	 	 else if (in == 2200) out = -2545;
	 	 	 else if (in == 2201) out = -2544;
	 	 	 else if (in == 2202) out = -2542;
	 	 	 else if (in == 2203) out = -2540;
	 	 	 else if (in == 2204) out = -2538;
	 	 	 else if (in == 2205) out = -2536;
	 	 	 else if (in == 2206) out = -2534;
	 	 	 else if (in == 2207) out = -2532;
	 	 	 else if (in == 2208) out = -2531;
	 	 	 else if (in == 2209) out = -2529;
	 	 	 else if (in == 2210) out = -2527;
	 	 	 else if (in == 2211) out = -2525;
	 	 	 else if (in == 2212) out = -2523;
	 	 	 else if (in == 2213) out = -2521;
	 	 	 else if (in == 2214) out = -2519;
	 	 	 else if (in == 2215) out = -2518;
	 	 	 else if (in == 2216) out = -2516;
	 	 	 else if (in == 2217) out = -2514;
	 	 	 else if (in == 2218) out = -2512;
	 	 	 else if (in == 2219) out = -2510;
	 	 	 else if (in == 2220) out = -2508;
	 	 	 else if (in == 2221) out = -2506;
	 	 	 else if (in == 2222) out = -2505;
	 	 	 else if (in == 2223) out = -2503;
	 	 	 else if (in == 2224) out = -2501;
	 	 	 else if (in == 2225) out = -2499;
	 	 	 else if (in == 2226) out = -2497;
	 	 	 else if (in == 2227) out = -2495;
	 	 	 else if (in == 2228) out = -2494;
	 	 	 else if (in == 2229) out = -2492;
	 	 	 else if (in == 2230) out = -2490;
	 	 	 else if (in == 2231) out = -2488;
	 	 	 else if (in == 2232) out = -2486;
	 	 	 else if (in == 2233) out = -2484;
	 	 	 else if (in == 2234) out = -2483;
	 	 	 else if (in == 2235) out = -2481;
	 	 	 else if (in == 2236) out = -2479;
	 	 	 else if (in == 2237) out = -2477;
	 	 	 else if (in == 2238) out = -2475;
	 	 	 else if (in == 2239) out = -2473;
	 	 	 else if (in == 2240) out = -2472;
	 	 	 else if (in == 2241) out = -2470;
	 	 	 else if (in == 2242) out = -2468;
	 	 	 else if (in == 2243) out = -2466;
	 	 	 else if (in == 2244) out = -2464;
	 	 	 else if (in == 2245) out = -2462;
	 	 	 else if (in == 2246) out = -2461;
	 	 	 else if (in == 2247) out = -2459;
	 	 	 else if (in == 2248) out = -2457;
	 	 	 else if (in == 2249) out = -2455;
	 	 	 else if (in == 2250) out = -2453;
	 	 	 else if (in == 2251) out = -2452;
	 	 	 else if (in == 2252) out = -2450;
	 	 	 else if (in == 2253) out = -2448;
	 	 	 else if (in == 2254) out = -2446;
	 	 	 else if (in == 2255) out = -2444;
	 	 	 else if (in == 2256) out = -2442;
	 	 	 else if (in == 2257) out = -2441;
	 	 	 else if (in == 2258) out = -2439;
	 	 	 else if (in == 2259) out = -2437;
	 	 	 else if (in == 2260) out = -2435;
	 	 	 else if (in == 2261) out = -2433;
	 	 	 else if (in == 2262) out = -2432;
	 	 	 else if (in == 2263) out = -2430;
	 	 	 else if (in == 2264) out = -2428;
	 	 	 else if (in == 2265) out = -2426;
	 	 	 else if (in == 2266) out = -2424;
	 	 	 else if (in == 2267) out = -2423;
	 	 	 else if (in == 2268) out = -2421;
	 	 	 else if (in == 2269) out = -2419;
	 	 	 else if (in == 2270) out = -2417;
	 	 	 else if (in == 2271) out = -2415;
	 	 	 else if (in == 2272) out = -2413;
	 	 	 else if (in == 2273) out = -2412;
	 	 	 else if (in == 2274) out = -2410;
	 	 	 else if (in == 2275) out = -2408;
	 	 	 else if (in == 2276) out = -2406;
	 	 	 else if (in == 2277) out = -2404;
	 	 	 else if (in == 2278) out = -2403;
	 	 	 else if (in == 2279) out = -2401;
	 	 	 else if (in == 2280) out = -2399;
	 	 	 else if (in == 2281) out = -2397;
	 	 	 else if (in == 2282) out = -2395;
	 	 	 else if (in == 2283) out = -2394;
	 	 	 else if (in == 2284) out = -2392;
	 	 	 else if (in == 2285) out = -2390;
	 	 	 else if (in == 2286) out = -2388;
	 	 	 else if (in == 2287) out = -2387;
	 	 	 else if (in == 2288) out = -2385;
	 	 	 else if (in == 2289) out = -2383;
	 	 	 else if (in == 2290) out = -2381;
	 	 	 else if (in == 2291) out = -2379;
	 	 	 else if (in == 2292) out = -2378;
	 	 	 else if (in == 2293) out = -2376;
	 	 	 else if (in == 2294) out = -2374;
	 	 	 else if (in == 2295) out = -2372;
	 	 	 else if (in == 2296) out = -2370;
	 	 	 else if (in == 2297) out = -2369;
	 	 	 else if (in == 2298) out = -2367;
	 	 	 else if (in == 2299) out = -2365;
	 	 	 else if (in == 2300) out = -2363;
	 	 	 else if (in == 2301) out = -2362;
	 	 	 else if (in == 2302) out = -2360;
	 	 	 else if (in == 2303) out = -2358;
	 	 	 else if (in == 2304) out = -2356;
	 	 	 else if (in == 2305) out = -2354;
	 	 	 else if (in == 2306) out = -2353;
	 	 	 else if (in == 2307) out = -2351;
	 	 	 else if (in == 2308) out = -2349;
	 	 	 else if (in == 2309) out = -2347;
	 	 	 else if (in == 2310) out = -2346;
	 	 	 else if (in == 2311) out = -2344;
	 	 	 else if (in == 2312) out = -2342;
	 	 	 else if (in == 2313) out = -2340;
	 	 	 else if (in == 2314) out = -2338;
	 	 	 else if (in == 2315) out = -2337;
	 	 	 else if (in == 2316) out = -2335;
	 	 	 else if (in == 2317) out = -2333;
	 	 	 else if (in == 2318) out = -2331;
	 	 	 else if (in == 2319) out = -2330;
	 	 	 else if (in == 2320) out = -2328;
	 	 	 else if (in == 2321) out = -2326;
	 	 	 else if (in == 2322) out = -2324;
	 	 	 else if (in == 2323) out = -2323;
	 	 	 else if (in == 2324) out = -2321;
	 	 	 else if (in == 2325) out = -2319;
	 	 	 else if (in == 2326) out = -2317;
	 	 	 else if (in == 2327) out = -2316;
	 	 	 else if (in == 2328) out = -2314;
	 	 	 else if (in == 2329) out = -2312;
	 	 	 else if (in == 2330) out = -2310;
	 	 	 else if (in == 2331) out = -2308;
	 	 	 else if (in == 2332) out = -2307;
	 	 	 else if (in == 2333) out = -2305;
	 	 	 else if (in == 2334) out = -2303;
	 	 	 else if (in == 2335) out = -2301;
	 	 	 else if (in == 2336) out = -2300;
	 	 	 else if (in == 2337) out = -2298;
	 	 	 else if (in == 2338) out = -2296;
	 	 	 else if (in == 2339) out = -2294;
	 	 	 else if (in == 2340) out = -2293;
	 	 	 else if (in == 2341) out = -2291;
	 	 	 else if (in == 2342) out = -2289;
	 	 	 else if (in == 2343) out = -2287;
	 	 	 else if (in == 2344) out = -2286;
	 	 	 else if (in == 2345) out = -2284;
	 	 	 else if (in == 2346) out = -2282;
	 	 	 else if (in == 2347) out = -2280;
	 	 	 else if (in == 2348) out = -2279;
	 	 	 else if (in == 2349) out = -2277;
	 	 	 else if (in == 2350) out = -2275;
	 	 	 else if (in == 2351) out = -2273;
	 	 	 else if (in == 2352) out = -2272;
	 	 	 else if (in == 2353) out = -2270;
	 	 	 else if (in == 2354) out = -2268;
	 	 	 else if (in == 2355) out = -2267;
	 	 	 else if (in == 2356) out = -2265;
	 	 	 else if (in == 2357) out = -2263;
	 	 	 else if (in == 2358) out = -2261;
	 	 	 else if (in == 2359) out = -2260;
	 	 	 else if (in == 2360) out = -2258;
	 	 	 else if (in == 2361) out = -2256;
	 	 	 else if (in == 2362) out = -2254;
	 	 	 else if (in == 2363) out = -2253;
	 	 	 else if (in == 2364) out = -2251;
	 	 	 else if (in == 2365) out = -2249;
	 	 	 else if (in == 2366) out = -2247;
	 	 	 else if (in == 2367) out = -2246;
	 	 	 else if (in == 2368) out = -2244;
	 	 	 else if (in == 2369) out = -2242;
	 	 	 else if (in == 2370) out = -2241;
	 	 	 else if (in == 2371) out = -2239;
	 	 	 else if (in == 2372) out = -2237;
	 	 	 else if (in == 2373) out = -2235;
	 	 	 else if (in == 2374) out = -2234;
	 	 	 else if (in == 2375) out = -2232;
	 	 	 else if (in == 2376) out = -2230;
	 	 	 else if (in == 2377) out = -2228;
	 	 	 else if (in == 2378) out = -2227;
	 	 	 else if (in == 2379) out = -2225;
	 	 	 else if (in == 2380) out = -2223;
	 	 	 else if (in == 2381) out = -2222;
	 	 	 else if (in == 2382) out = -2220;
	 	 	 else if (in == 2383) out = -2218;
	 	 	 else if (in == 2384) out = -2216;
	 	 	 else if (in == 2385) out = -2215;
	 	 	 else if (in == 2386) out = -2213;
	 	 	 else if (in == 2387) out = -2211;
	 	 	 else if (in == 2388) out = -2210;
	 	 	 else if (in == 2389) out = -2208;
	 	 	 else if (in == 2390) out = -2206;
	 	 	 else if (in == 2391) out = -2204;
	 	 	 else if (in == 2392) out = -2203;
	 	 	 else if (in == 2393) out = -2201;
	 	 	 else if (in == 2394) out = -2199;
	 	 	 else if (in == 2395) out = -2198;
	 	 	 else if (in == 2396) out = -2196;
	 	 	 else if (in == 2397) out = -2194;
	 	 	 else if (in == 2398) out = -2192;
	 	 	 else if (in == 2399) out = -2191;
	 	 	 else if (in == 2400) out = -2189;
	 	 	 else if (in == 2401) out = -2187;
	 	 	 else if (in == 2402) out = -2186;
	 	 	 else if (in == 2403) out = -2184;
	 	 	 else if (in == 2404) out = -2182;
	 	 	 else if (in == 2405) out = -2180;
	 	 	 else if (in == 2406) out = -2179;
	 	 	 else if (in == 2407) out = -2177;
	 	 	 else if (in == 2408) out = -2175;
	 	 	 else if (in == 2409) out = -2174;
	 	 	 else if (in == 2410) out = -2172;
	 	 	 else if (in == 2411) out = -2170;
	 	 	 else if (in == 2412) out = -2169;
	 	 	 else if (in == 2413) out = -2167;
	 	 	 else if (in == 2414) out = -2165;
	 	 	 else if (in == 2415) out = -2163;
	 	 	 else if (in == 2416) out = -2162;
	 	 	 else if (in == 2417) out = -2160;
	 	 	 else if (in == 2418) out = -2158;
	 	 	 else if (in == 2419) out = -2157;
	 	 	 else if (in == 2420) out = -2155;
	 	 	 else if (in == 2421) out = -2153;
	 	 	 else if (in == 2422) out = -2152;
	 	 	 else if (in == 2423) out = -2150;
	 	 	 else if (in == 2424) out = -2148;
	 	 	 else if (in == 2425) out = -2147;
	 	 	 else if (in == 2426) out = -2145;
	 	 	 else if (in == 2427) out = -2143;
	 	 	 else if (in == 2428) out = -2141;
	 	 	 else if (in == 2429) out = -2140;
	 	 	 else if (in == 2430) out = -2138;
	 	 	 else if (in == 2431) out = -2136;
	 	 	 else if (in == 2432) out = -2135;
	 	 	 else if (in == 2433) out = -2133;
	 	 	 else if (in == 2434) out = -2131;
	 	 	 else if (in == 2435) out = -2130;
	 	 	 else if (in == 2436) out = -2128;
	 	 	 else if (in == 2437) out = -2126;
	 	 	 else if (in == 2438) out = -2125;
	 	 	 else if (in == 2439) out = -2123;
	 	 	 else if (in == 2440) out = -2121;
	 	 	 else if (in == 2441) out = -2120;
	 	 	 else if (in == 2442) out = -2118;
	 	 	 else if (in == 2443) out = -2116;
	 	 	 else if (in == 2444) out = -2115;
	 	 	 else if (in == 2445) out = -2113;
	 	 	 else if (in == 2446) out = -2111;
	 	 	 else if (in == 2447) out = -2110;
	 	 	 else if (in == 2448) out = -2108;
	 	 	 else if (in == 2449) out = -2106;
	 	 	 else if (in == 2450) out = -2105;
	 	 	 else if (in == 2451) out = -2103;
	 	 	 else if (in == 2452) out = -2101;
	 	 	 else if (in == 2453) out = -2100;
	 	 	 else if (in == 2454) out = -2098;
	 	 	 else if (in == 2455) out = -2096;
	 	 	 else if (in == 2456) out = -2095;
	 	 	 else if (in == 2457) out = -2093;
	 	 	 else if (in == 2458) out = -2091;
	 	 	 else if (in == 2459) out = -2090;
	 	 	 else if (in == 2460) out = -2088;
	 	 	 else if (in == 2461) out = -2086;
	 	 	 else if (in == 2462) out = -2085;
	 	 	 else if (in == 2463) out = -2083;
	 	 	 else if (in == 2464) out = -2081;
	 	 	 else if (in == 2465) out = -2080;
	 	 	 else if (in == 2466) out = -2078;
	 	 	 else if (in == 2467) out = -2076;
	 	 	 else if (in == 2468) out = -2075;
	 	 	 else if (in == 2469) out = -2073;
	 	 	 else if (in == 2470) out = -2071;
	 	 	 else if (in == 2471) out = -2070;
	 	 	 else if (in == 2472) out = -2068;
	 	 	 else if (in == 2473) out = -2066;
	 	 	 else if (in == 2474) out = -2065;
	 	 	 else if (in == 2475) out = -2063;
	 	 	 else if (in == 2476) out = -2061;
	 	 	 else if (in == 2477) out = -2060;
	 	 	 else if (in == 2478) out = -2058;
	 	 	 else if (in == 2479) out = -2056;
	 	 	 else if (in == 2480) out = -2055;
	 	 	 else if (in == 2481) out = -2053;
	 	 	 else if (in == 2482) out = -2051;
	 	 	 else if (in == 2483) out = -2050;
	 	 	 else if (in == 2484) out = -2048;
	 	 	 else if (in == 2485) out = -2046;
	 	 	 else if (in == 2486) out = -2045;
	 	 	 else if (in == 2487) out = -2043;
	 	 	 else if (in == 2488) out = -2041;
	 	 	 else if (in == 2489) out = -2040;
	 	 	 else if (in == 2490) out = -2038;
	 	 	 else if (in == 2491) out = -2037;
	 	 	 else if (in == 2492) out = -2035;
	 	 	 else if (in == 2493) out = -2033;
	 	 	 else if (in == 2494) out = -2032;
	 	 	 else if (in == 2495) out = -2030;
	 	 	 else if (in == 2496) out = -2028;
	 	 	 else if (in == 2497) out = -2027;
	 	 	 else if (in == 2498) out = -2025;
	 	 	 else if (in == 2499) out = -2023;
	 	 	 else if (in == 2500) out = -2022;
	 	 	 else if (in == 2501) out = -2020;
	 	 	 else if (in == 2502) out = -2019;
	 	 	 else if (in == 2503) out = -2017;
	 	 	 else if (in == 2504) out = -2015;
	 	 	 else if (in == 2505) out = -2014;
	 	 	 else if (in == 2506) out = -2012;
	 	 	 else if (in == 2507) out = -2010;
	 	 	 else if (in == 2508) out = -2009;
	 	 	 else if (in == 2509) out = -2007;
	 	 	 else if (in == 2510) out = -2005;
	 	 	 else if (in == 2511) out = -2004;
	 	 	 else if (in == 2512) out = -2002;
	 	 	 else if (in == 2513) out = -2001;
	 	 	 else if (in == 2514) out = -1999;
	 	 	 else if (in == 2515) out = -1997;
	 	 	 else if (in == 2516) out = -1996;
	 	 	 else if (in == 2517) out = -1994;
	 	 	 else if (in == 2518) out = -1992;
	 	 	 else if (in == 2519) out = -1991;
	 	 	 else if (in == 2520) out = -1989;
	 	 	 else if (in == 2521) out = -1988;
	 	 	 else if (in == 2522) out = -1986;
	 	 	 else if (in == 2523) out = -1984;
	 	 	 else if (in == 2524) out = -1983;
	 	 	 else if (in == 2525) out = -1981;
	 	 	 else if (in == 2526) out = -1979;
	 	 	 else if (in == 2527) out = -1978;
	 	 	 else if (in == 2528) out = -1976;
	 	 	 else if (in == 2529) out = -1975;
	 	 	 else if (in == 2530) out = -1973;
	 	 	 else if (in == 2531) out = -1971;
	 	 	 else if (in == 2532) out = -1970;
	 	 	 else if (in == 2533) out = -1968;
	 	 	 else if (in == 2534) out = -1966;
	 	 	 else if (in == 2535) out = -1965;
	 	 	 else if (in == 2536) out = -1963;
	 	 	 else if (in == 2537) out = -1962;
	 	 	 else if (in == 2538) out = -1960;
	 	 	 else if (in == 2539) out = -1958;
	 	 	 else if (in == 2540) out = -1957;
	 	 	 else if (in == 2541) out = -1955;
	 	 	 else if (in == 2542) out = -1954;
	 	 	 else if (in == 2543) out = -1952;
	 	 	 else if (in == 2544) out = -1950;
	 	 	 else if (in == 2545) out = -1949;
	 	 	 else if (in == 2546) out = -1947;
	 	 	 else if (in == 2547) out = -1945;
	 	 	 else if (in == 2548) out = -1944;
	 	 	 else if (in == 2549) out = -1942;
	 	 	 else if (in == 2550) out = -1941;
	 	 	 else if (in == 2551) out = -1939;
	 	 	 else if (in == 2552) out = -1937;
	 	 	 else if (in == 2553) out = -1936;
	 	 	 else if (in == 2554) out = -1934;
	 	 	 else if (in == 2555) out = -1933;
	 	 	 else if (in == 2556) out = -1931;
	 	 	 else if (in == 2557) out = -1929;
	 	 	 else if (in == 2558) out = -1928;
	 	 	 else if (in == 2559) out = -1926;
	 	 	 else if (in == 2560) out = -1925;
	 	 	 else if (in == 2561) out = -1923;
	 	 	 else if (in == 2562) out = -1921;
	 	 	 else if (in == 2563) out = -1920;
	 	 	 else if (in == 2564) out = -1918;
	 	 	 else if (in == 2565) out = -1917;
	 	 	 else if (in == 2566) out = -1915;
	 	 	 else if (in == 2567) out = -1913;
	 	 	 else if (in == 2568) out = -1912;
	 	 	 else if (in == 2569) out = -1910;
	 	 	 else if (in == 2570) out = -1909;
	 	 	 else if (in == 2571) out = -1907;
	 	 	 else if (in == 2572) out = -1905;
	 	 	 else if (in == 2573) out = -1904;
	 	 	 else if (in == 2574) out = -1902;
	 	 	 else if (in == 2575) out = -1901;
	 	 	 else if (in == 2576) out = -1899;
	 	 	 else if (in == 2577) out = -1898;
	 	 	 else if (in == 2578) out = -1896;
	 	 	 else if (in == 2579) out = -1894;
	 	 	 else if (in == 2580) out = -1893;
	 	 	 else if (in == 2581) out = -1891;
	 	 	 else if (in == 2582) out = -1890;
	 	 	 else if (in == 2583) out = -1888;
	 	 	 else if (in == 2584) out = -1886;
	 	 	 else if (in == 2585) out = -1885;
	 	 	 else if (in == 2586) out = -1883;
	 	 	 else if (in == 2587) out = -1882;
	 	 	 else if (in == 2588) out = -1880;
	 	 	 else if (in == 2589) out = -1878;
	 	 	 else if (in == 2590) out = -1877;
	 	 	 else if (in == 2591) out = -1875;
	 	 	 else if (in == 2592) out = -1874;
	 	 	 else if (in == 2593) out = -1872;
	 	 	 else if (in == 2594) out = -1871;
	 	 	 else if (in == 2595) out = -1869;
	 	 	 else if (in == 2596) out = -1867;
	 	 	 else if (in == 2597) out = -1866;
	 	 	 else if (in == 2598) out = -1864;
	 	 	 else if (in == 2599) out = -1863;
	 	 	 else if (in == 2600) out = -1861;
	 	 	 else if (in == 2601) out = -1860;
	 	 	 else if (in == 2602) out = -1858;
	 	 	 else if (in == 2603) out = -1856;
	 	 	 else if (in == 2604) out = -1855;
	 	 	 else if (in == 2605) out = -1853;
	 	 	 else if (in == 2606) out = -1852;
	 	 	 else if (in == 2607) out = -1850;
	 	 	 else if (in == 2608) out = -1849;
	 	 	 else if (in == 2609) out = -1847;
	 	 	 else if (in == 2610) out = -1845;
	 	 	 else if (in == 2611) out = -1844;
	 	 	 else if (in == 2612) out = -1842;
	 	 	 else if (in == 2613) out = -1841;
	 	 	 else if (in == 2614) out = -1839;
	 	 	 else if (in == 2615) out = -1838;
	 	 	 else if (in == 2616) out = -1836;
	 	 	 else if (in == 2617) out = -1834;
	 	 	 else if (in == 2618) out = -1833;
	 	 	 else if (in == 2619) out = -1831;
	 	 	 else if (in == 2620) out = -1830;
	 	 	 else if (in == 2621) out = -1828;
	 	 	 else if (in == 2622) out = -1827;
	 	 	 else if (in == 2623) out = -1825;
	 	 	 else if (in == 2624) out = -1823;
	 	 	 else if (in == 2625) out = -1822;
	 	 	 else if (in == 2626) out = -1820;
	 	 	 else if (in == 2627) out = -1819;
	 	 	 else if (in == 2628) out = -1817;
	 	 	 else if (in == 2629) out = -1816;
	 	 	 else if (in == 2630) out = -1814;
	 	 	 else if (in == 2631) out = -1813;
	 	 	 else if (in == 2632) out = -1811;
	 	 	 else if (in == 2633) out = -1809;
	 	 	 else if (in == 2634) out = -1808;
	 	 	 else if (in == 2635) out = -1806;
	 	 	 else if (in == 2636) out = -1805;
	 	 	 else if (in == 2637) out = -1803;
	 	 	 else if (in == 2638) out = -1802;
	 	 	 else if (in == 2639) out = -1800;
	 	 	 else if (in == 2640) out = -1799;
	 	 	 else if (in == 2641) out = -1797;
	 	 	 else if (in == 2642) out = -1795;
	 	 	 else if (in == 2643) out = -1794;
	 	 	 else if (in == 2644) out = -1792;
	 	 	 else if (in == 2645) out = -1791;
	 	 	 else if (in == 2646) out = -1789;
	 	 	 else if (in == 2647) out = -1788;
	 	 	 else if (in == 2648) out = -1786;
	 	 	 else if (in == 2649) out = -1785;
	 	 	 else if (in == 2650) out = -1783;
	 	 	 else if (in == 2651) out = -1782;
	 	 	 else if (in == 2652) out = -1780;
	 	 	 else if (in == 2653) out = -1778;
	 	 	 else if (in == 2654) out = -1777;
	 	 	 else if (in == 2655) out = -1775;
	 	 	 else if (in == 2656) out = -1774;
	 	 	 else if (in == 2657) out = -1772;
	 	 	 else if (in == 2658) out = -1771;
	 	 	 else if (in == 2659) out = -1769;
	 	 	 else if (in == 2660) out = -1768;
	 	 	 else if (in == 2661) out = -1766;
	 	 	 else if (in == 2662) out = -1765;
	 	 	 else if (in == 2663) out = -1763;
	 	 	 else if (in == 2664) out = -1762;
	 	 	 else if (in == 2665) out = -1760;
	 	 	 else if (in == 2666) out = -1758;
	 	 	 else if (in == 2667) out = -1757;
	 	 	 else if (in == 2668) out = -1755;
	 	 	 else if (in == 2669) out = -1754;
	 	 	 else if (in == 2670) out = -1752;
	 	 	 else if (in == 2671) out = -1751;
	 	 	 else if (in == 2672) out = -1749;
	 	 	 else if (in == 2673) out = -1748;
	 	 	 else if (in == 2674) out = -1746;
	 	 	 else if (in == 2675) out = -1745;
	 	 	 else if (in == 2676) out = -1743;
	 	 	 else if (in == 2677) out = -1742;
	 	 	 else if (in == 2678) out = -1740;
	 	 	 else if (in == 2679) out = -1739;
	 	 	 else if (in == 2680) out = -1737;
	 	 	 else if (in == 2681) out = -1735;
	 	 	 else if (in == 2682) out = -1734;
	 	 	 else if (in == 2683) out = -1732;
	 	 	 else if (in == 2684) out = -1731;
	 	 	 else if (in == 2685) out = -1729;
	 	 	 else if (in == 2686) out = -1728;
	 	 	 else if (in == 2687) out = -1726;
	 	 	 else if (in == 2688) out = -1725;
	 	 	 else if (in == 2689) out = -1723;
	 	 	 else if (in == 2690) out = -1722;
	 	 	 else if (in == 2691) out = -1720;
	 	 	 else if (in == 2692) out = -1719;
	 	 	 else if (in == 2693) out = -1717;
	 	 	 else if (in == 2694) out = -1716;
	 	 	 else if (in == 2695) out = -1714;
	 	 	 else if (in == 2696) out = -1713;
	 	 	 else if (in == 2697) out = -1711;
	 	 	 else if (in == 2698) out = -1710;
	 	 	 else if (in == 2699) out = -1708;
	 	 	 else if (in == 2700) out = -1707;
	 	 	 else if (in == 2701) out = -1705;
	 	 	 else if (in == 2702) out = -1704;
	 	 	 else if (in == 2703) out = -1702;
	 	 	 else if (in == 2704) out = -1700;
	 	 	 else if (in == 2705) out = -1699;
	 	 	 else if (in == 2706) out = -1697;
	 	 	 else if (in == 2707) out = -1696;
	 	 	 else if (in == 2708) out = -1694;
	 	 	 else if (in == 2709) out = -1693;
	 	 	 else if (in == 2710) out = -1691;
	 	 	 else if (in == 2711) out = -1690;
	 	 	 else if (in == 2712) out = -1688;
	 	 	 else if (in == 2713) out = -1687;
	 	 	 else if (in == 2714) out = -1685;
	 	 	 else if (in == 2715) out = -1684;
	 	 	 else if (in == 2716) out = -1682;
	 	 	 else if (in == 2717) out = -1681;
	 	 	 else if (in == 2718) out = -1679;
	 	 	 else if (in == 2719) out = -1678;
	 	 	 else if (in == 2720) out = -1676;
	 	 	 else if (in == 2721) out = -1675;
	 	 	 else if (in == 2722) out = -1673;
	 	 	 else if (in == 2723) out = -1672;
	 	 	 else if (in == 2724) out = -1670;
	 	 	 else if (in == 2725) out = -1669;
	 	 	 else if (in == 2726) out = -1667;
	 	 	 else if (in == 2727) out = -1666;
	 	 	 else if (in == 2728) out = -1664;
	 	 	 else if (in == 2729) out = -1663;
	 	 	 else if (in == 2730) out = -1661;
	 	 	 else if (in == 2731) out = -1660;
	 	 	 else if (in == 2732) out = -1658;
	 	 	 else if (in == 2733) out = -1657;
	 	 	 else if (in == 2734) out = -1655;
	 	 	 else if (in == 2735) out = -1654;
	 	 	 else if (in == 2736) out = -1652;
	 	 	 else if (in == 2737) out = -1651;
	 	 	 else if (in == 2738) out = -1649;
	 	 	 else if (in == 2739) out = -1648;
	 	 	 else if (in == 2740) out = -1646;
	 	 	 else if (in == 2741) out = -1645;
	 	 	 else if (in == 2742) out = -1643;
	 	 	 else if (in == 2743) out = -1642;
	 	 	 else if (in == 2744) out = -1640;
	 	 	 else if (in == 2745) out = -1639;
	 	 	 else if (in == 2746) out = -1637;
	 	 	 else if (in == 2747) out = -1636;
	 	 	 else if (in == 2748) out = -1634;
	 	 	 else if (in == 2749) out = -1633;
	 	 	 else if (in == 2750) out = -1631;
	 	 	 else if (in == 2751) out = -1630;
	 	 	 else if (in == 2752) out = -1628;
	 	 	 else if (in == 2753) out = -1627;
	 	 	 else if (in == 2754) out = -1625;
	 	 	 else if (in == 2755) out = -1624;
	 	 	 else if (in == 2756) out = -1622;
	 	 	 else if (in == 2757) out = -1621;
	 	 	 else if (in == 2758) out = -1619;
	 	 	 else if (in == 2759) out = -1618;
	 	 	 else if (in == 2760) out = -1617;
	 	 	 else if (in == 2761) out = -1615;
	 	 	 else if (in == 2762) out = -1614;
	 	 	 else if (in == 2763) out = -1612;
	 	 	 else if (in == 2764) out = -1611;
	 	 	 else if (in == 2765) out = -1609;
	 	 	 else if (in == 2766) out = -1608;
	 	 	 else if (in == 2767) out = -1606;
	 	 	 else if (in == 2768) out = -1605;
	 	 	 else if (in == 2769) out = -1603;
	 	 	 else if (in == 2770) out = -1602;
	 	 	 else if (in == 2771) out = -1600;
	 	 	 else if (in == 2772) out = -1599;
	 	 	 else if (in == 2773) out = -1597;
	 	 	 else if (in == 2774) out = -1596;
	 	 	 else if (in == 2775) out = -1594;
	 	 	 else if (in == 2776) out = -1593;
	 	 	 else if (in == 2777) out = -1591;
	 	 	 else if (in == 2778) out = -1590;
	 	 	 else if (in == 2779) out = -1588;
	 	 	 else if (in == 2780) out = -1587;
	 	 	 else if (in == 2781) out = -1585;
	 	 	 else if (in == 2782) out = -1584;
	 	 	 else if (in == 2783) out = -1583;
	 	 	 else if (in == 2784) out = -1581;
	 	 	 else if (in == 2785) out = -1580;
	 	 	 else if (in == 2786) out = -1578;
	 	 	 else if (in == 2787) out = -1577;
	 	 	 else if (in == 2788) out = -1575;
	 	 	 else if (in == 2789) out = -1574;
	 	 	 else if (in == 2790) out = -1572;
	 	 	 else if (in == 2791) out = -1571;
	 	 	 else if (in == 2792) out = -1569;
	 	 	 else if (in == 2793) out = -1568;
	 	 	 else if (in == 2794) out = -1566;
	 	 	 else if (in == 2795) out = -1565;
	 	 	 else if (in == 2796) out = -1563;
	 	 	 else if (in == 2797) out = -1562;
	 	 	 else if (in == 2798) out = -1561;
	 	 	 else if (in == 2799) out = -1559;
	 	 	 else if (in == 2800) out = -1558;
	 	 	 else if (in == 2801) out = -1556;
	 	 	 else if (in == 2802) out = -1555;
	 	 	 else if (in == 2803) out = -1553;
	 	 	 else if (in == 2804) out = -1552;
	 	 	 else if (in == 2805) out = -1550;
	 	 	 else if (in == 2806) out = -1549;
	 	 	 else if (in == 2807) out = -1547;
	 	 	 else if (in == 2808) out = -1546;
	 	 	 else if (in == 2809) out = -1544;
	 	 	 else if (in == 2810) out = -1543;
	 	 	 else if (in == 2811) out = -1542;
	 	 	 else if (in == 2812) out = -1540;
	 	 	 else if (in == 2813) out = -1539;
	 	 	 else if (in == 2814) out = -1537;
	 	 	 else if (in == 2815) out = -1536;
	 	 	 else if (in == 2816) out = -1534;
	 	 	 else if (in == 2817) out = -1533;
	 	 	 else if (in == 2818) out = -1531;
	 	 	 else if (in == 2819) out = -1530;
	 	 	 else if (in == 2820) out = -1528;
	 	 	 else if (in == 2821) out = -1527;
	 	 	 else if (in == 2822) out = -1526;
	 	 	 else if (in == 2823) out = -1524;
	 	 	 else if (in == 2824) out = -1523;
	 	 	 else if (in == 2825) out = -1521;
	 	 	 else if (in == 2826) out = -1520;
	 	 	 else if (in == 2827) out = -1518;
	 	 	 else if (in == 2828) out = -1517;
	 	 	 else if (in == 2829) out = -1515;
	 	 	 else if (in == 2830) out = -1514;
	 	 	 else if (in == 2831) out = -1512;
	 	 	 else if (in == 2832) out = -1511;
	 	 	 else if (in == 2833) out = -1510;
	 	 	 else if (in == 2834) out = -1508;
	 	 	 else if (in == 2835) out = -1507;
	 	 	 else if (in == 2836) out = -1505;
	 	 	 else if (in == 2837) out = -1504;
	 	 	 else if (in == 2838) out = -1502;
	 	 	 else if (in == 2839) out = -1501;
	 	 	 else if (in == 2840) out = -1499;
	 	 	 else if (in == 2841) out = -1498;
	 	 	 else if (in == 2842) out = -1497;
	 	 	 else if (in == 2843) out = -1495;
	 	 	 else if (in == 2844) out = -1494;
	 	 	 else if (in == 2845) out = -1492;
	 	 	 else if (in == 2846) out = -1491;
	 	 	 else if (in == 2847) out = -1489;
	 	 	 else if (in == 2848) out = -1488;
	 	 	 else if (in == 2849) out = -1487;
	 	 	 else if (in == 2850) out = -1485;
	 	 	 else if (in == 2851) out = -1484;
	 	 	 else if (in == 2852) out = -1482;
	 	 	 else if (in == 2853) out = -1481;
	 	 	 else if (in == 2854) out = -1479;
	 	 	 else if (in == 2855) out = -1478;
	 	 	 else if (in == 2856) out = -1476;
	 	 	 else if (in == 2857) out = -1475;
	 	 	 else if (in == 2858) out = -1474;
	 	 	 else if (in == 2859) out = -1472;
	 	 	 else if (in == 2860) out = -1471;
	 	 	 else if (in == 2861) out = -1469;
	 	 	 else if (in == 2862) out = -1468;
	 	 	 else if (in == 2863) out = -1466;
	 	 	 else if (in == 2864) out = -1465;
	 	 	 else if (in == 2865) out = -1464;
	 	 	 else if (in == 2866) out = -1462;
	 	 	 else if (in == 2867) out = -1461;
	 	 	 else if (in == 2868) out = -1459;
	 	 	 else if (in == 2869) out = -1458;
	 	 	 else if (in == 2870) out = -1456;
	 	 	 else if (in == 2871) out = -1455;
	 	 	 else if (in == 2872) out = -1454;
	 	 	 else if (in == 2873) out = -1452;
	 	 	 else if (in == 2874) out = -1451;
	 	 	 else if (in == 2875) out = -1449;
	 	 	 else if (in == 2876) out = -1448;
	 	 	 else if (in == 2877) out = -1446;
	 	 	 else if (in == 2878) out = -1445;
	 	 	 else if (in == 2879) out = -1444;
	 	 	 else if (in == 2880) out = -1442;
	 	 	 else if (in == 2881) out = -1441;
	 	 	 else if (in == 2882) out = -1439;
	 	 	 else if (in == 2883) out = -1438;
	 	 	 else if (in == 2884) out = -1437;
	 	 	 else if (in == 2885) out = -1435;
	 	 	 else if (in == 2886) out = -1434;
	 	 	 else if (in == 2887) out = -1432;
	 	 	 else if (in == 2888) out = -1431;
	 	 	 else if (in == 2889) out = -1429;
	 	 	 else if (in == 2890) out = -1428;
	 	 	 else if (in == 2891) out = -1427;
	 	 	 else if (in == 2892) out = -1425;
	 	 	 else if (in == 2893) out = -1424;
	 	 	 else if (in == 2894) out = -1422;
	 	 	 else if (in == 2895) out = -1421;
	 	 	 else if (in == 2896) out = -1420;
	 	 	 else if (in == 2897) out = -1418;
	 	 	 else if (in == 2898) out = -1417;
	 	 	 else if (in == 2899) out = -1415;
	 	 	 else if (in == 2900) out = -1414;
	 	 	 else if (in == 2901) out = -1412;
	 	 	 else if (in == 2902) out = -1411;
	 	 	 else if (in == 2903) out = -1410;
	 	 	 else if (in == 2904) out = -1408;
	 	 	 else if (in == 2905) out = -1407;
	 	 	 else if (in == 2906) out = -1405;
	 	 	 else if (in == 2907) out = -1404;
	 	 	 else if (in == 2908) out = -1403;
	 	 	 else if (in == 2909) out = -1401;
	 	 	 else if (in == 2910) out = -1400;
	 	 	 else if (in == 2911) out = -1398;
	 	 	 else if (in == 2912) out = -1397;
	 	 	 else if (in == 2913) out = -1396;
	 	 	 else if (in == 2914) out = -1394;
	 	 	 else if (in == 2915) out = -1393;
	 	 	 else if (in == 2916) out = -1391;
	 	 	 else if (in == 2917) out = -1390;
	 	 	 else if (in == 2918) out = -1389;
	 	 	 else if (in == 2919) out = -1387;
	 	 	 else if (in == 2920) out = -1386;
	 	 	 else if (in == 2921) out = -1384;
	 	 	 else if (in == 2922) out = -1383;
	 	 	 else if (in == 2923) out = -1381;
	 	 	 else if (in == 2924) out = -1380;
	 	 	 else if (in == 2925) out = -1379;
	 	 	 else if (in == 2926) out = -1377;
	 	 	 else if (in == 2927) out = -1376;
	 	 	 else if (in == 2928) out = -1374;
	 	 	 else if (in == 2929) out = -1373;
	 	 	 else if (in == 2930) out = -1372;
	 	 	 else if (in == 2931) out = -1370;
	 	 	 else if (in == 2932) out = -1369;
	 	 	 else if (in == 2933) out = -1368;
	 	 	 else if (in == 2934) out = -1366;
	 	 	 else if (in == 2935) out = -1365;
	 	 	 else if (in == 2936) out = -1363;
	 	 	 else if (in == 2937) out = -1362;
	 	 	 else if (in == 2938) out = -1361;
	 	 	 else if (in == 2939) out = -1359;
	 	 	 else if (in == 2940) out = -1358;
	 	 	 else if (in == 2941) out = -1356;
	 	 	 else if (in == 2942) out = -1355;
	 	 	 else if (in == 2943) out = -1354;
	 	 	 else if (in == 2944) out = -1352;
	 	 	 else if (in == 2945) out = -1351;
	 	 	 else if (in == 2946) out = -1349;
	 	 	 else if (in == 2947) out = -1348;
	 	 	 else if (in == 2948) out = -1347;
	 	 	 else if (in == 2949) out = -1345;
	 	 	 else if (in == 2950) out = -1344;
	 	 	 else if (in == 2951) out = -1342;
	 	 	 else if (in == 2952) out = -1341;
	 	 	 else if (in == 2953) out = -1340;
	 	 	 else if (in == 2954) out = -1338;
	 	 	 else if (in == 2955) out = -1337;
	 	 	 else if (in == 2956) out = -1336;
	 	 	 else if (in == 2957) out = -1334;
	 	 	 else if (in == 2958) out = -1333;
	 	 	 else if (in == 2959) out = -1331;
	 	 	 else if (in == 2960) out = -1330;
	 	 	 else if (in == 2961) out = -1329;
	 	 	 else if (in == 2962) out = -1327;
	 	 	 else if (in == 2963) out = -1326;
	 	 	 else if (in == 2964) out = -1324;
	 	 	 else if (in == 2965) out = -1323;
	 	 	 else if (in == 2966) out = -1322;
	 	 	 else if (in == 2967) out = -1320;
	 	 	 else if (in == 2968) out = -1319;
	 	 	 else if (in == 2969) out = -1318;
	 	 	 else if (in == 2970) out = -1316;
	 	 	 else if (in == 2971) out = -1315;
	 	 	 else if (in == 2972) out = -1313;
	 	 	 else if (in == 2973) out = -1312;
	 	 	 else if (in == 2974) out = -1311;
	 	 	 else if (in == 2975) out = -1309;
	 	 	 else if (in == 2976) out = -1308;
	 	 	 else if (in == 2977) out = -1307;
	 	 	 else if (in == 2978) out = -1305;
	 	 	 else if (in == 2979) out = -1304;
	 	 	 else if (in == 2980) out = -1302;
	 	 	 else if (in == 2981) out = -1301;
	 	 	 else if (in == 2982) out = -1300;
	 	 	 else if (in == 2983) out = -1298;
	 	 	 else if (in == 2984) out = -1297;
	 	 	 else if (in == 2985) out = -1296;
	 	 	 else if (in == 2986) out = -1294;
	 	 	 else if (in == 2987) out = -1293;
	 	 	 else if (in == 2988) out = -1291;
	 	 	 else if (in == 2989) out = -1290;
	 	 	 else if (in == 2990) out = -1289;
	 	 	 else if (in == 2991) out = -1287;
	 	 	 else if (in == 2992) out = -1286;
	 	 	 else if (in == 2993) out = -1285;
	 	 	 else if (in == 2994) out = -1283;
	 	 	 else if (in == 2995) out = -1282;
	 	 	 else if (in == 2996) out = -1280;
	 	 	 else if (in == 2997) out = -1279;
	 	 	 else if (in == 2998) out = -1278;
	 	 	 else if (in == 2999) out = -1276;
	 	 	 else if (in == 3000) out = -1275;
	 	 	 else if (in == 3001) out = -1274;
	 	 	 else if (in == 3002) out = -1272;
	 	 	 else if (in == 3003) out = -1271;
	 	 	 else if (in == 3004) out = -1270;
	 	 	 else if (in == 3005) out = -1268;
	 	 	 else if (in == 3006) out = -1267;
	 	 	 else if (in == 3007) out = -1265;
	 	 	 else if (in == 3008) out = -1264;
	 	 	 else if (in == 3009) out = -1263;
	 	 	 else if (in == 3010) out = -1261;
	 	 	 else if (in == 3011) out = -1260;
	 	 	 else if (in == 3012) out = -1259;
	 	 	 else if (in == 3013) out = -1257;
	 	 	 else if (in == 3014) out = -1256;
	 	 	 else if (in == 3015) out = -1255;
	 	 	 else if (in == 3016) out = -1253;
	 	 	 else if (in == 3017) out = -1252;
	 	 	 else if (in == 3018) out = -1250;
	 	 	 else if (in == 3019) out = -1249;
	 	 	 else if (in == 3020) out = -1248;
	 	 	 else if (in == 3021) out = -1246;
	 	 	 else if (in == 3022) out = -1245;
	 	 	 else if (in == 3023) out = -1244;
	 	 	 else if (in == 3024) out = -1242;
	 	 	 else if (in == 3025) out = -1241;
	 	 	 else if (in == 3026) out = -1240;
	 	 	 else if (in == 3027) out = -1238;
	 	 	 else if (in == 3028) out = -1237;
	 	 	 else if (in == 3029) out = -1236;
	 	 	 else if (in == 3030) out = -1234;
	 	 	 else if (in == 3031) out = -1233;
	 	 	 else if (in == 3032) out = -1232;
	 	 	 else if (in == 3033) out = -1230;
	 	 	 else if (in == 3034) out = -1229;
	 	 	 else if (in == 3035) out = -1227;
	 	 	 else if (in == 3036) out = -1226;
	 	 	 else if (in == 3037) out = -1225;
	 	 	 else if (in == 3038) out = -1223;
	 	 	 else if (in == 3039) out = -1222;
	 	 	 else if (in == 3040) out = -1221;
	 	 	 else if (in == 3041) out = -1219;
	 	 	 else if (in == 3042) out = -1218;
	 	 	 else if (in == 3043) out = -1217;
	 	 	 else if (in == 3044) out = -1215;
	 	 	 else if (in == 3045) out = -1214;
	 	 	 else if (in == 3046) out = -1213;
	 	 	 else if (in == 3047) out = -1211;
	 	 	 else if (in == 3048) out = -1210;
	 	 	 else if (in == 3049) out = -1209;
	 	 	 else if (in == 3050) out = -1207;
	 	 	 else if (in == 3051) out = -1206;
	 	 	 else if (in == 3052) out = -1205;
	 	 	 else if (in == 3053) out = -1203;
	 	 	 else if (in == 3054) out = -1202;
	 	 	 else if (in == 3055) out = -1201;
	 	 	 else if (in == 3056) out = -1199;
	 	 	 else if (in == 3057) out = -1198;
	 	 	 else if (in == 3058) out = -1197;
	 	 	 else if (in == 3059) out = -1195;
	 	 	 else if (in == 3060) out = -1194;
	 	 	 else if (in == 3061) out = -1193;
	 	 	 else if (in == 3062) out = -1191;
	 	 	 else if (in == 3063) out = -1190;
	 	 	 else if (in == 3064) out = -1189;
	 	 	 else if (in == 3065) out = -1187;
	 	 	 else if (in == 3066) out = -1186;
	 	 	 else if (in == 3067) out = -1185;
	 	 	 else if (in == 3068) out = -1183;
	 	 	 else if (in == 3069) out = -1182;
	 	 	 else if (in == 3070) out = -1181;
	 	 	 else if (in == 3071) out = -1179;
	 	 	 else if (in == 3072) out = -1178;
	 	 	 else if (in == 3073) out = -1177;
	 	 	 else if (in == 3074) out = -1175;
	 	 	 else if (in == 3075) out = -1174;
	 	 	 else if (in == 3076) out = -1173;
	 	 	 else if (in == 3077) out = -1171;
	 	 	 else if (in == 3078) out = -1170;
	 	 	 else if (in == 3079) out = -1169;
	 	 	 else if (in == 3080) out = -1167;
	 	 	 else if (in == 3081) out = -1166;
	 	 	 else if (in == 3082) out = -1165;
	 	 	 else if (in == 3083) out = -1163;
	 	 	 else if (in == 3084) out = -1162;
	 	 	 else if (in == 3085) out = -1161;
	 	 	 else if (in == 3086) out = -1159;
	 	 	 else if (in == 3087) out = -1158;
	 	 	 else if (in == 3088) out = -1157;
	 	 	 else if (in == 3089) out = -1155;
	 	 	 else if (in == 3090) out = -1154;
	 	 	 else if (in == 3091) out = -1153;
	 	 	 else if (in == 3092) out = -1151;
	 	 	 else if (in == 3093) out = -1150;
	 	 	 else if (in == 3094) out = -1149;
	 	 	 else if (in == 3095) out = -1147;
	 	 	 else if (in == 3096) out = -1146;
	 	 	 else if (in == 3097) out = -1145;
	 	 	 else if (in == 3098) out = -1143;
	 	 	 else if (in == 3099) out = -1142;
	 	 	 else if (in == 3100) out = -1141;
	 	 	 else if (in == 3101) out = -1139;
	 	 	 else if (in == 3102) out = -1138;
	 	 	 else if (in == 3103) out = -1137;
	 	 	 else if (in == 3104) out = -1135;
	 	 	 else if (in == 3105) out = -1134;
	 	 	 else if (in == 3106) out = -1133;
	 	 	 else if (in == 3107) out = -1131;
	 	 	 else if (in == 3108) out = -1130;
	 	 	 else if (in == 3109) out = -1129;
	 	 	 else if (in == 3110) out = -1127;
	 	 	 else if (in == 3111) out = -1126;
	 	 	 else if (in == 3112) out = -1125;
	 	 	 else if (in == 3113) out = -1124;
	 	 	 else if (in == 3114) out = -1122;
	 	 	 else if (in == 3115) out = -1121;
	 	 	 else if (in == 3116) out = -1120;
	 	 	 else if (in == 3117) out = -1118;
	 	 	 else if (in == 3118) out = -1117;
	 	 	 else if (in == 3119) out = -1116;
	 	 	 else if (in == 3120) out = -1114;
	 	 	 else if (in == 3121) out = -1113;
	 	 	 else if (in == 3122) out = -1112;
	 	 	 else if (in == 3123) out = -1110;
	 	 	 else if (in == 3124) out = -1109;
	 	 	 else if (in == 3125) out = -1108;
	 	 	 else if (in == 3126) out = -1106;
	 	 	 else if (in == 3127) out = -1105;
	 	 	 else if (in == 3128) out = -1104;
	 	 	 else if (in == 3129) out = -1103;
	 	 	 else if (in == 3130) out = -1101;
	 	 	 else if (in == 3131) out = -1100;
	 	 	 else if (in == 3132) out = -1099;
	 	 	 else if (in == 3133) out = -1097;
	 	 	 else if (in == 3134) out = -1096;
	 	 	 else if (in == 3135) out = -1095;
	 	 	 else if (in == 3136) out = -1093;
	 	 	 else if (in == 3137) out = -1092;
	 	 	 else if (in == 3138) out = -1091;
	 	 	 else if (in == 3139) out = -1089;
	 	 	 else if (in == 3140) out = -1088;
	 	 	 else if (in == 3141) out = -1087;
	 	 	 else if (in == 3142) out = -1086;
	 	 	 else if (in == 3143) out = -1084;
	 	 	 else if (in == 3144) out = -1083;
	 	 	 else if (in == 3145) out = -1082;
	 	 	 else if (in == 3146) out = -1080;
	 	 	 else if (in == 3147) out = -1079;
	 	 	 else if (in == 3148) out = -1078;
	 	 	 else if (in == 3149) out = -1076;
	 	 	 else if (in == 3150) out = -1075;
	 	 	 else if (in == 3151) out = -1074;
	 	 	 else if (in == 3152) out = -1073;
	 	 	 else if (in == 3153) out = -1071;
	 	 	 else if (in == 3154) out = -1070;
	 	 	 else if (in == 3155) out = -1069;
	 	 	 else if (in == 3156) out = -1067;
	 	 	 else if (in == 3157) out = -1066;
	 	 	 else if (in == 3158) out = -1065;
	 	 	 else if (in == 3159) out = -1063;
	 	 	 else if (in == 3160) out = -1062;
	 	 	 else if (in == 3161) out = -1061;
	 	 	 else if (in == 3162) out = -1060;
	 	 	 else if (in == 3163) out = -1058;
	 	 	 else if (in == 3164) out = -1057;
	 	 	 else if (in == 3165) out = -1056;
	 	 	 else if (in == 3166) out = -1054;
	 	 	 else if (in == 3167) out = -1053;
	 	 	 else if (in == 3168) out = -1052;
	 	 	 else if (in == 3169) out = -1051;
	 	 	 else if (in == 3170) out = -1049;
	 	 	 else if (in == 3171) out = -1048;
	 	 	 else if (in == 3172) out = -1047;
	 	 	 else if (in == 3173) out = -1045;
	 	 	 else if (in == 3174) out = -1044;
	 	 	 else if (in == 3175) out = -1043;
	 	 	 else if (in == 3176) out = -1041;
	 	 	 else if (in == 3177) out = -1040;
	 	 	 else if (in == 3178) out = -1039;
	 	 	 else if (in == 3179) out = -1038;
	 	 	 else if (in == 3180) out = -1036;
	 	 	 else if (in == 3181) out = -1035;
	 	 	 else if (in == 3182) out = -1034;
	 	 	 else if (in == 3183) out = -1032;
	 	 	 else if (in == 3184) out = -1031;
	 	 	 else if (in == 3185) out = -1030;
	 	 	 else if (in == 3186) out = -1029;
	 	 	 else if (in == 3187) out = -1027;
	 	 	 else if (in == 3188) out = -1026;
	 	 	 else if (in == 3189) out = -1025;
	 	 	 else if (in == 3190) out = -1023;
	 	 	 else if (in == 3191) out = -1022;
	 	 	 else if (in == 3192) out = -1021;
	 	 	 else if (in == 3193) out = -1020;
	 	 	 else if (in == 3194) out = -1018;
	 	 	 else if (in == 3195) out = -1017;
	 	 	 else if (in == 3196) out = -1016;
	 	 	 else if (in == 3197) out = -1014;
	 	 	 else if (in == 3198) out = -1013;
	 	 	 else if (in == 3199) out = -1012;
	 	 	 else if (in == 3200) out = -1011;
	 	 	 else if (in == 3201) out = -1009;
	 	 	 else if (in == 3202) out = -1008;
	 	 	 else if (in == 3203) out = -1007;
	 	 	 else if (in == 3204) out = -1006;
	 	 	 else if (in == 3205) out = -1004;
	 	 	 else if (in == 3206) out = -1003;
	 	 	 else if (in == 3207) out = -1002;
	 	 	 else if (in == 3208) out = -1000;
	 	 	 else if (in == 3209) out = -999;
	 	 	 else if (in == 3210) out = -998;
	 	 	 else if (in == 3211) out = -997;
	 	 	 else if (in == 3212) out = -995;
	 	 	 else if (in == 3213) out = -994;
	 	 	 else if (in == 3214) out = -993;
	 	 	 else if (in == 3215) out = -991;
	 	 	 else if (in == 3216) out = -990;
	 	 	 else if (in == 3217) out = -989;
	 	 	 else if (in == 3218) out = -988;
	 	 	 else if (in == 3219) out = -986;
	 	 	 else if (in == 3220) out = -985;
	 	 	 else if (in == 3221) out = -984;
	 	 	 else if (in == 3222) out = -983;
	 	 	 else if (in == 3223) out = -981;
	 	 	 else if (in == 3224) out = -980;
	 	 	 else if (in == 3225) out = -979;
	 	 	 else if (in == 3226) out = -977;
	 	 	 else if (in == 3227) out = -976;
	 	 	 else if (in == 3228) out = -975;
	 	 	 else if (in == 3229) out = -974;
	 	 	 else if (in == 3230) out = -972;
	 	 	 else if (in == 3231) out = -971;
	 	 	 else if (in == 3232) out = -970;
	 	 	 else if (in == 3233) out = -969;
	 	 	 else if (in == 3234) out = -967;
	 	 	 else if (in == 3235) out = -966;
	 	 	 else if (in == 3236) out = -965;
	 	 	 else if (in == 3237) out = -964;
	 	 	 else if (in == 3238) out = -962;
	 	 	 else if (in == 3239) out = -961;
	 	 	 else if (in == 3240) out = -960;
	 	 	 else if (in == 3241) out = -958;
	 	 	 else if (in == 3242) out = -957;
	 	 	 else if (in == 3243) out = -956;
	 	 	 else if (in == 3244) out = -955;
	 	 	 else if (in == 3245) out = -953;
	 	 	 else if (in == 3246) out = -952;
	 	 	 else if (in == 3247) out = -951;
	 	 	 else if (in == 3248) out = -950;
	 	 	 else if (in == 3249) out = -948;
	 	 	 else if (in == 3250) out = -947;
	 	 	 else if (in == 3251) out = -946;
	 	 	 else if (in == 3252) out = -945;
	 	 	 else if (in == 3253) out = -943;
	 	 	 else if (in == 3254) out = -942;
	 	 	 else if (in == 3255) out = -941;
	 	 	 else if (in == 3256) out = -940;
	 	 	 else if (in == 3257) out = -938;
	 	 	 else if (in == 3258) out = -937;
	 	 	 else if (in == 3259) out = -936;
	 	 	 else if (in == 3260) out = -935;
	 	 	 else if (in == 3261) out = -933;
	 	 	 else if (in == 3262) out = -932;
	 	 	 else if (in == 3263) out = -931;
	 	 	 else if (in == 3264) out = -930;
	 	 	 else if (in == 3265) out = -928;
	 	 	 else if (in == 3266) out = -927;
	 	 	 else if (in == 3267) out = -926;
	 	 	 else if (in == 3268) out = -925;
	 	 	 else if (in == 3269) out = -923;
	 	 	 else if (in == 3270) out = -922;
	 	 	 else if (in == 3271) out = -921;
	 	 	 else if (in == 3272) out = -920;
	 	 	 else if (in == 3273) out = -918;
	 	 	 else if (in == 3274) out = -917;
	 	 	 else if (in == 3275) out = -916;
	 	 	 else if (in == 3276) out = -914;
	 	 	 else if (in == 3277) out = -913;
	 	 	 else if (in == 3278) out = -912;
	 	 	 else if (in == 3279) out = -911;
	 	 	 else if (in == 3280) out = -909;
	 	 	 else if (in == 3281) out = -908;
	 	 	 else if (in == 3282) out = -907;
	 	 	 else if (in == 3283) out = -906;
	 	 	 else if (in == 3284) out = -905;
	 	 	 else if (in == 3285) out = -903;
	 	 	 else if (in == 3286) out = -902;
	 	 	 else if (in == 3287) out = -901;
	 	 	 else if (in == 3288) out = -900;
	 	 	 else if (in == 3289) out = -898;
	 	 	 else if (in == 3290) out = -897;
	 	 	 else if (in == 3291) out = -896;
	 	 	 else if (in == 3292) out = -895;
	 	 	 else if (in == 3293) out = -893;
	 	 	 else if (in == 3294) out = -892;
	 	 	 else if (in == 3295) out = -891;
	 	 	 else if (in == 3296) out = -890;
	 	 	 else if (in == 3297) out = -888;
	 	 	 else if (in == 3298) out = -887;
	 	 	 else if (in == 3299) out = -886;
	 	 	 else if (in == 3300) out = -885;
	 	 	 else if (in == 3301) out = -883;
	 	 	 else if (in == 3302) out = -882;
	 	 	 else if (in == 3303) out = -881;
	 	 	 else if (in == 3304) out = -880;
	 	 	 else if (in == 3305) out = -878;
	 	 	 else if (in == 3306) out = -877;
	 	 	 else if (in == 3307) out = -876;
	 	 	 else if (in == 3308) out = -875;
	 	 	 else if (in == 3309) out = -873;
	 	 	 else if (in == 3310) out = -872;
	 	 	 else if (in == 3311) out = -871;
	 	 	 else if (in == 3312) out = -870;
	 	 	 else if (in == 3313) out = -868;
	 	 	 else if (in == 3314) out = -867;
	 	 	 else if (in == 3315) out = -866;
	 	 	 else if (in == 3316) out = -865;
	 	 	 else if (in == 3317) out = -864;
	 	 	 else if (in == 3318) out = -862;
	 	 	 else if (in == 3319) out = -861;
	 	 	 else if (in == 3320) out = -860;
	 	 	 else if (in == 3321) out = -859;
	 	 	 else if (in == 3322) out = -857;
	 	 	 else if (in == 3323) out = -856;
	 	 	 else if (in == 3324) out = -855;
	 	 	 else if (in == 3325) out = -854;
	 	 	 else if (in == 3326) out = -852;
	 	 	 else if (in == 3327) out = -851;
	 	 	 else if (in == 3328) out = -850;
	 	 	 else if (in == 3329) out = -849;
	 	 	 else if (in == 3330) out = -848;
	 	 	 else if (in == 3331) out = -846;
	 	 	 else if (in == 3332) out = -845;
	 	 	 else if (in == 3333) out = -844;
	 	 	 else if (in == 3334) out = -843;
	 	 	 else if (in == 3335) out = -841;
	 	 	 else if (in == 3336) out = -840;
	 	 	 else if (in == 3337) out = -839;
	 	 	 else if (in == 3338) out = -838;
	 	 	 else if (in == 3339) out = -836;
	 	 	 else if (in == 3340) out = -835;
	 	 	 else if (in == 3341) out = -834;
	 	 	 else if (in == 3342) out = -833;
	 	 	 else if (in == 3343) out = -832;
	 	 	 else if (in == 3344) out = -830;
	 	 	 else if (in == 3345) out = -829;
	 	 	 else if (in == 3346) out = -828;
	 	 	 else if (in == 3347) out = -827;
	 	 	 else if (in == 3348) out = -825;
	 	 	 else if (in == 3349) out = -824;
	 	 	 else if (in == 3350) out = -823;
	 	 	 else if (in == 3351) out = -822;
	 	 	 else if (in == 3352) out = -821;
	 	 	 else if (in == 3353) out = -819;
	 	 	 else if (in == 3354) out = -818;
	 	 	 else if (in == 3355) out = -817;
	 	 	 else if (in == 3356) out = -816;
	 	 	 else if (in == 3357) out = -814;
	 	 	 else if (in == 3358) out = -813;
	 	 	 else if (in == 3359) out = -812;
	 	 	 else if (in == 3360) out = -811;
	 	 	 else if (in == 3361) out = -810;
	 	 	 else if (in == 3362) out = -808;
	 	 	 else if (in == 3363) out = -807;
	 	 	 else if (in == 3364) out = -806;
	 	 	 else if (in == 3365) out = -805;
	 	 	 else if (in == 3366) out = -803;
	 	 	 else if (in == 3367) out = -802;
	 	 	 else if (in == 3368) out = -801;
	 	 	 else if (in == 3369) out = -800;
	 	 	 else if (in == 3370) out = -799;
	 	 	 else if (in == 3371) out = -797;
	 	 	 else if (in == 3372) out = -796;
	 	 	 else if (in == 3373) out = -795;
	 	 	 else if (in == 3374) out = -794;
	 	 	 else if (in == 3375) out = -793;
	 	 	 else if (in == 3376) out = -791;
	 	 	 else if (in == 3377) out = -790;
	 	 	 else if (in == 3378) out = -789;
	 	 	 else if (in == 3379) out = -788;
	 	 	 else if (in == 3380) out = -786;
	 	 	 else if (in == 3381) out = -785;
	 	 	 else if (in == 3382) out = -784;
	 	 	 else if (in == 3383) out = -783;
	 	 	 else if (in == 3384) out = -782;
	 	 	 else if (in == 3385) out = -780;
	 	 	 else if (in == 3386) out = -779;
	 	 	 else if (in == 3387) out = -778;
	 	 	 else if (in == 3388) out = -777;
	 	 	 else if (in == 3389) out = -776;
	 	 	 else if (in == 3390) out = -774;
	 	 	 else if (in == 3391) out = -773;
	 	 	 else if (in == 3392) out = -772;
	 	 	 else if (in == 3393) out = -771;
	 	 	 else if (in == 3394) out = -770;
	 	 	 else if (in == 3395) out = -768;
	 	 	 else if (in == 3396) out = -767;
	 	 	 else if (in == 3397) out = -766;
	 	 	 else if (in == 3398) out = -765;
	 	 	 else if (in == 3399) out = -764;
	 	 	 else if (in == 3400) out = -762;
	 	 	 else if (in == 3401) out = -761;
	 	 	 else if (in == 3402) out = -760;
	 	 	 else if (in == 3403) out = -759;
	 	 	 else if (in == 3404) out = -758;
	 	 	 else if (in == 3405) out = -756;
	 	 	 else if (in == 3406) out = -755;
	 	 	 else if (in == 3407) out = -754;
	 	 	 else if (in == 3408) out = -753;
	 	 	 else if (in == 3409) out = -751;
	 	 	 else if (in == 3410) out = -750;
	 	 	 else if (in == 3411) out = -749;
	 	 	 else if (in == 3412) out = -748;
	 	 	 else if (in == 3413) out = -747;
	 	 	 else if (in == 3414) out = -745;
	 	 	 else if (in == 3415) out = -744;
	 	 	 else if (in == 3416) out = -743;
	 	 	 else if (in == 3417) out = -742;
	 	 	 else if (in == 3418) out = -741;
	 	 	 else if (in == 3419) out = -739;
	 	 	 else if (in == 3420) out = -738;
	 	 	 else if (in == 3421) out = -737;
	 	 	 else if (in == 3422) out = -736;
	 	 	 else if (in == 3423) out = -735;
	 	 	 else if (in == 3424) out = -734;
	 	 	 else if (in == 3425) out = -732;
	 	 	 else if (in == 3426) out = -731;
	 	 	 else if (in == 3427) out = -730;
	 	 	 else if (in == 3428) out = -729;
	 	 	 else if (in == 3429) out = -728;
	 	 	 else if (in == 3430) out = -726;
	 	 	 else if (in == 3431) out = -725;
	 	 	 else if (in == 3432) out = -724;
	 	 	 else if (in == 3433) out = -723;
	 	 	 else if (in == 3434) out = -722;
	 	 	 else if (in == 3435) out = -720;
	 	 	 else if (in == 3436) out = -719;
	 	 	 else if (in == 3437) out = -718;
	 	 	 else if (in == 3438) out = -717;
	 	 	 else if (in == 3439) out = -716;
	 	 	 else if (in == 3440) out = -714;
	 	 	 else if (in == 3441) out = -713;
	 	 	 else if (in == 3442) out = -712;
	 	 	 else if (in == 3443) out = -711;
	 	 	 else if (in == 3444) out = -710;
	 	 	 else if (in == 3445) out = -708;
	 	 	 else if (in == 3446) out = -707;
	 	 	 else if (in == 3447) out = -706;
	 	 	 else if (in == 3448) out = -705;
	 	 	 else if (in == 3449) out = -704;
	 	 	 else if (in == 3450) out = -703;
	 	 	 else if (in == 3451) out = -701;
	 	 	 else if (in == 3452) out = -700;
	 	 	 else if (in == 3453) out = -699;
	 	 	 else if (in == 3454) out = -698;
	 	 	 else if (in == 3455) out = -697;
	 	 	 else if (in == 3456) out = -695;
	 	 	 else if (in == 3457) out = -694;
	 	 	 else if (in == 3458) out = -693;
	 	 	 else if (in == 3459) out = -692;
	 	 	 else if (in == 3460) out = -691;
	 	 	 else if (in == 3461) out = -689;
	 	 	 else if (in == 3462) out = -688;
	 	 	 else if (in == 3463) out = -687;
	 	 	 else if (in == 3464) out = -686;
	 	 	 else if (in == 3465) out = -685;
	 	 	 else if (in == 3466) out = -684;
	 	 	 else if (in == 3467) out = -682;
	 	 	 else if (in == 3468) out = -681;
	 	 	 else if (in == 3469) out = -680;
	 	 	 else if (in == 3470) out = -679;
	 	 	 else if (in == 3471) out = -678;
	 	 	 else if (in == 3472) out = -676;
	 	 	 else if (in == 3473) out = -675;
	 	 	 else if (in == 3474) out = -674;
	 	 	 else if (in == 3475) out = -673;
	 	 	 else if (in == 3476) out = -672;
	 	 	 else if (in == 3477) out = -671;
	 	 	 else if (in == 3478) out = -669;
	 	 	 else if (in == 3479) out = -668;
	 	 	 else if (in == 3480) out = -667;
	 	 	 else if (in == 3481) out = -666;
	 	 	 else if (in == 3482) out = -665;
	 	 	 else if (in == 3483) out = -664;
	 	 	 else if (in == 3484) out = -662;
	 	 	 else if (in == 3485) out = -661;
	 	 	 else if (in == 3486) out = -660;
	 	 	 else if (in == 3487) out = -659;
	 	 	 else if (in == 3488) out = -658;
	 	 	 else if (in == 3489) out = -656;
	 	 	 else if (in == 3490) out = -655;
	 	 	 else if (in == 3491) out = -654;
	 	 	 else if (in == 3492) out = -653;
	 	 	 else if (in == 3493) out = -652;
	 	 	 else if (in == 3494) out = -651;
	 	 	 else if (in == 3495) out = -649;
	 	 	 else if (in == 3496) out = -648;
	 	 	 else if (in == 3497) out = -647;
	 	 	 else if (in == 3498) out = -646;
	 	 	 else if (in == 3499) out = -645;
	 	 	 else if (in == 3500) out = -644;
	 	 	 else if (in == 3501) out = -642;
	 	 	 else if (in == 3502) out = -641;
	 	 	 else if (in == 3503) out = -640;
	 	 	 else if (in == 3504) out = -639;
	 	 	 else if (in == 3505) out = -638;
	 	 	 else if (in == 3506) out = -637;
	 	 	 else if (in == 3507) out = -635;
	 	 	 else if (in == 3508) out = -634;
	 	 	 else if (in == 3509) out = -633;
	 	 	 else if (in == 3510) out = -632;
	 	 	 else if (in == 3511) out = -631;
	 	 	 else if (in == 3512) out = -630;
	 	 	 else if (in == 3513) out = -628;
	 	 	 else if (in == 3514) out = -627;
	 	 	 else if (in == 3515) out = -626;
	 	 	 else if (in == 3516) out = -625;
	 	 	 else if (in == 3517) out = -624;
	 	 	 else if (in == 3518) out = -623;
	 	 	 else if (in == 3519) out = -621;
	 	 	 else if (in == 3520) out = -620;
	 	 	 else if (in == 3521) out = -619;
	 	 	 else if (in == 3522) out = -618;
	 	 	 else if (in == 3523) out = -617;
	 	 	 else if (in == 3524) out = -616;
	 	 	 else if (in == 3525) out = -614;
	 	 	 else if (in == 3526) out = -613;
	 	 	 else if (in == 3527) out = -612;
	 	 	 else if (in == 3528) out = -611;
	 	 	 else if (in == 3529) out = -610;
	 	 	 else if (in == 3530) out = -609;
	 	 	 else if (in == 3531) out = -607;
	 	 	 else if (in == 3532) out = -606;
	 	 	 else if (in == 3533) out = -605;
	 	 	 else if (in == 3534) out = -604;
	 	 	 else if (in == 3535) out = -603;
	 	 	 else if (in == 3536) out = -602;
	 	 	 else if (in == 3537) out = -601;
	 	 	 else if (in == 3538) out = -599;
	 	 	 else if (in == 3539) out = -598;
	 	 	 else if (in == 3540) out = -597;
	 	 	 else if (in == 3541) out = -596;
	 	 	 else if (in == 3542) out = -595;
	 	 	 else if (in == 3543) out = -594;
	 	 	 else if (in == 3544) out = -592;
	 	 	 else if (in == 3545) out = -591;
	 	 	 else if (in == 3546) out = -590;
	 	 	 else if (in == 3547) out = -589;
	 	 	 else if (in == 3548) out = -588;
	 	 	 else if (in == 3549) out = -587;
	 	 	 else if (in == 3550) out = -585;
	 	 	 else if (in == 3551) out = -584;
	 	 	 else if (in == 3552) out = -583;
	 	 	 else if (in == 3553) out = -582;
	 	 	 else if (in == 3554) out = -581;
	 	 	 else if (in == 3555) out = -580;
	 	 	 else if (in == 3556) out = -579;
	 	 	 else if (in == 3557) out = -577;
	 	 	 else if (in == 3558) out = -576;
	 	 	 else if (in == 3559) out = -575;
	 	 	 else if (in == 3560) out = -574;
	 	 	 else if (in == 3561) out = -573;
	 	 	 else if (in == 3562) out = -572;
	 	 	 else if (in == 3563) out = -571;
	 	 	 else if (in == 3564) out = -569;
	 	 	 else if (in == 3565) out = -568;
	 	 	 else if (in == 3566) out = -567;
	 	 	 else if (in == 3567) out = -566;
	 	 	 else if (in == 3568) out = -565;
	 	 	 else if (in == 3569) out = -564;
	 	 	 else if (in == 3570) out = -562;
	 	 	 else if (in == 3571) out = -561;
	 	 	 else if (in == 3572) out = -560;
	 	 	 else if (in == 3573) out = -559;
	 	 	 else if (in == 3574) out = -558;
	 	 	 else if (in == 3575) out = -557;
	 	 	 else if (in == 3576) out = -556;
	 	 	 else if (in == 3577) out = -554;
	 	 	 else if (in == 3578) out = -553;
	 	 	 else if (in == 3579) out = -552;
	 	 	 else if (in == 3580) out = -551;
	 	 	 else if (in == 3581) out = -550;
	 	 	 else if (in == 3582) out = -549;
	 	 	 else if (in == 3583) out = -548;
	 	 	 else if (in == 3584) out = -546;
	 	 	 else if (in == 3585) out = -545;
	 	 	 else if (in == 3586) out = -544;
	 	 	 else if (in == 3587) out = -543;
	 	 	 else if (in == 3588) out = -542;
	 	 	 else if (in == 3589) out = -541;
	 	 	 else if (in == 3590) out = -540;
	 	 	 else if (in == 3591) out = -538;
	 	 	 else if (in == 3592) out = -537;
	 	 	 else if (in == 3593) out = -536;
	 	 	 else if (in == 3594) out = -535;
	 	 	 else if (in == 3595) out = -534;
	 	 	 else if (in == 3596) out = -533;
	 	 	 else if (in == 3597) out = -532;
	 	 	 else if (in == 3598) out = -530;
	 	 	 else if (in == 3599) out = -529;
	 	 	 else if (in == 3600) out = -528;
	 	 	 else if (in == 3601) out = -527;
	 	 	 else if (in == 3602) out = -526;
	 	 	 else if (in == 3603) out = -525;
	 	 	 else if (in == 3604) out = -524;
	 	 	 else if (in == 3605) out = -523;
	 	 	 else if (in == 3606) out = -521;
	 	 	 else if (in == 3607) out = -520;
	 	 	 else if (in == 3608) out = -519;
	 	 	 else if (in == 3609) out = -518;
	 	 	 else if (in == 3610) out = -517;
	 	 	 else if (in == 3611) out = -516;
	 	 	 else if (in == 3612) out = -515;
	 	 	 else if (in == 3613) out = -513;
	 	 	 else if (in == 3614) out = -512;
	 	 	 else if (in == 3615) out = -511;
	 	 	 else if (in == 3616) out = -510;
	 	 	 else if (in == 3617) out = -509;
	 	 	 else if (in == 3618) out = -508;
	 	 	 else if (in == 3619) out = -507;
	 	 	 else if (in == 3620) out = -506;
	 	 	 else if (in == 3621) out = -504;
	 	 	 else if (in == 3622) out = -503;
	 	 	 else if (in == 3623) out = -502;
	 	 	 else if (in == 3624) out = -501;
	 	 	 else if (in == 3625) out = -500;
	 	 	 else if (in == 3626) out = -499;
	 	 	 else if (in == 3627) out = -498;
	 	 	 else if (in == 3628) out = -496;
	 	 	 else if (in == 3629) out = -495;
	 	 	 else if (in == 3630) out = -494;
	 	 	 else if (in == 3631) out = -493;
	 	 	 else if (in == 3632) out = -492;
	 	 	 else if (in == 3633) out = -491;
	 	 	 else if (in == 3634) out = -490;
	 	 	 else if (in == 3635) out = -489;
	 	 	 else if (in == 3636) out = -487;
	 	 	 else if (in == 3637) out = -486;
	 	 	 else if (in == 3638) out = -485;
	 	 	 else if (in == 3639) out = -484;
	 	 	 else if (in == 3640) out = -483;
	 	 	 else if (in == 3641) out = -482;
	 	 	 else if (in == 3642) out = -481;
	 	 	 else if (in == 3643) out = -480;
	 	 	 else if (in == 3644) out = -478;
	 	 	 else if (in == 3645) out = -477;
	 	 	 else if (in == 3646) out = -476;
	 	 	 else if (in == 3647) out = -475;
	 	 	 else if (in == 3648) out = -474;
	 	 	 else if (in == 3649) out = -473;
	 	 	 else if (in == 3650) out = -472;
	 	 	 else if (in == 3651) out = -471;
	 	 	 else if (in == 3652) out = -469;
	 	 	 else if (in == 3653) out = -468;
	 	 	 else if (in == 3654) out = -467;
	 	 	 else if (in == 3655) out = -466;
	 	 	 else if (in == 3656) out = -465;
	 	 	 else if (in == 3657) out = -464;
	 	 	 else if (in == 3658) out = -463;
	 	 	 else if (in == 3659) out = -462;
	 	 	 else if (in == 3660) out = -460;
	 	 	 else if (in == 3661) out = -459;
	 	 	 else if (in == 3662) out = -458;
	 	 	 else if (in == 3663) out = -457;
	 	 	 else if (in == 3664) out = -456;
	 	 	 else if (in == 3665) out = -455;
	 	 	 else if (in == 3666) out = -454;
	 	 	 else if (in == 3667) out = -453;
	 	 	 else if (in == 3668) out = -452;
	 	 	 else if (in == 3669) out = -450;
	 	 	 else if (in == 3670) out = -449;
	 	 	 else if (in == 3671) out = -448;
	 	 	 else if (in == 3672) out = -447;
	 	 	 else if (in == 3673) out = -446;
	 	 	 else if (in == 3674) out = -445;
	 	 	 else if (in == 3675) out = -444;
	 	 	 else if (in == 3676) out = -443;
	 	 	 else if (in == 3677) out = -442;
	 	 	 else if (in == 3678) out = -440;
	 	 	 else if (in == 3679) out = -439;
	 	 	 else if (in == 3680) out = -438;
	 	 	 else if (in == 3681) out = -437;
	 	 	 else if (in == 3682) out = -436;
	 	 	 else if (in == 3683) out = -435;
	 	 	 else if (in == 3684) out = -434;
	 	 	 else if (in == 3685) out = -433;
	 	 	 else if (in == 3686) out = -432;
	 	 	 else if (in == 3687) out = -430;
	 	 	 else if (in == 3688) out = -429;
	 	 	 else if (in == 3689) out = -428;
	 	 	 else if (in == 3690) out = -427;
	 	 	 else if (in == 3691) out = -426;
	 	 	 else if (in == 3692) out = -425;
	 	 	 else if (in == 3693) out = -424;
	 	 	 else if (in == 3694) out = -423;
	 	 	 else if (in == 3695) out = -422;
	 	 	 else if (in == 3696) out = -420;
	 	 	 else if (in == 3697) out = -419;
	 	 	 else if (in == 3698) out = -418;
	 	 	 else if (in == 3699) out = -417;
	 	 	 else if (in == 3700) out = -416;
	 	 	 else if (in == 3701) out = -415;
	 	 	 else if (in == 3702) out = -414;
	 	 	 else if (in == 3703) out = -413;
	 	 	 else if (in == 3704) out = -412;
	 	 	 else if (in == 3705) out = -410;
	 	 	 else if (in == 3706) out = -409;
	 	 	 else if (in == 3707) out = -408;
	 	 	 else if (in == 3708) out = -407;
	 	 	 else if (in == 3709) out = -406;
	 	 	 else if (in == 3710) out = -405;
	 	 	 else if (in == 3711) out = -404;
	 	 	 else if (in == 3712) out = -403;
	 	 	 else if (in == 3713) out = -402;
	 	 	 else if (in == 3714) out = -401;
	 	 	 else if (in == 3715) out = -399;
	 	 	 else if (in == 3716) out = -398;
	 	 	 else if (in == 3717) out = -397;
	 	 	 else if (in == 3718) out = -396;
	 	 	 else if (in == 3719) out = -395;
	 	 	 else if (in == 3720) out = -394;
	 	 	 else if (in == 3721) out = -393;
	 	 	 else if (in == 3722) out = -392;
	 	 	 else if (in == 3723) out = -391;
	 	 	 else if (in == 3724) out = -389;
	 	 	 else if (in == 3725) out = -388;
	 	 	 else if (in == 3726) out = -387;
	 	 	 else if (in == 3727) out = -386;
	 	 	 else if (in == 3728) out = -385;
	 	 	 else if (in == 3729) out = -384;
	 	 	 else if (in == 3730) out = -383;
	 	 	 else if (in == 3731) out = -382;
	 	 	 else if (in == 3732) out = -381;
	 	 	 else if (in == 3733) out = -380;
	 	 	 else if (in == 3734) out = -379;
	 	 	 else if (in == 3735) out = -377;
	 	 	 else if (in == 3736) out = -376;
	 	 	 else if (in == 3737) out = -375;
	 	 	 else if (in == 3738) out = -374;
	 	 	 else if (in == 3739) out = -373;
	 	 	 else if (in == 3740) out = -372;
	 	 	 else if (in == 3741) out = -371;
	 	 	 else if (in == 3742) out = -370;
	 	 	 else if (in == 3743) out = -369;
	 	 	 else if (in == 3744) out = -368;
	 	 	 else if (in == 3745) out = -366;
	 	 	 else if (in == 3746) out = -365;
	 	 	 else if (in == 3747) out = -364;
	 	 	 else if (in == 3748) out = -363;
	 	 	 else if (in == 3749) out = -362;
	 	 	 else if (in == 3750) out = -361;
	 	 	 else if (in == 3751) out = -360;
	 	 	 else if (in == 3752) out = -359;
	 	 	 else if (in == 3753) out = -358;
	 	 	 else if (in == 3754) out = -357;
	 	 	 else if (in == 3755) out = -356;
	 	 	 else if (in == 3756) out = -354;
	 	 	 else if (in == 3757) out = -353;
	 	 	 else if (in == 3758) out = -352;
	 	 	 else if (in == 3759) out = -351;
	 	 	 else if (in == 3760) out = -350;
	 	 	 else if (in == 3761) out = -349;
	 	 	 else if (in == 3762) out = -348;
	 	 	 else if (in == 3763) out = -347;
	 	 	 else if (in == 3764) out = -346;
	 	 	 else if (in == 3765) out = -345;
	 	 	 else if (in == 3766) out = -344;
	 	 	 else if (in == 3767) out = -342;
	 	 	 else if (in == 3768) out = -341;
	 	 	 else if (in == 3769) out = -340;
	 	 	 else if (in == 3770) out = -339;
	 	 	 else if (in == 3771) out = -338;
	 	 	 else if (in == 3772) out = -337;
	 	 	 else if (in == 3773) out = -336;
	 	 	 else if (in == 3774) out = -335;
	 	 	 else if (in == 3775) out = -334;
	 	 	 else if (in == 3776) out = -333;
	 	 	 else if (in == 3777) out = -332;
	 	 	 else if (in == 3778) out = -331;
	 	 	 else if (in == 3779) out = -329;
	 	 	 else if (in == 3780) out = -328;
	 	 	 else if (in == 3781) out = -327;
	 	 	 else if (in == 3782) out = -326;
	 	 	 else if (in == 3783) out = -325;
	 	 	 else if (in == 3784) out = -324;
	 	 	 else if (in == 3785) out = -323;
	 	 	 else if (in == 3786) out = -322;
	 	 	 else if (in == 3787) out = -321;
	 	 	 else if (in == 3788) out = -320;
	 	 	 else if (in == 3789) out = -319;
	 	 	 else if (in == 3790) out = -318;
	 	 	 else if (in == 3791) out = -316;
	 	 	 else if (in == 3792) out = -315;
	 	 	 else if (in == 3793) out = -314;
	 	 	 else if (in == 3794) out = -313;
	 	 	 else if (in == 3795) out = -312;
	 	 	 else if (in == 3796) out = -311;
	 	 	 else if (in == 3797) out = -310;
	 	 	 else if (in == 3798) out = -309;
	 	 	 else if (in == 3799) out = -308;
	 	 	 else if (in == 3800) out = -307;
	 	 	 else if (in == 3801) out = -306;
	 	 	 else if (in == 3802) out = -305;
	 	 	 else if (in == 3803) out = -304;
	 	 	 else if (in == 3804) out = -302;
	 	 	 else if (in == 3805) out = -301;
	 	 	 else if (in == 3806) out = -300;
	 	 	 else if (in == 3807) out = -299;
	 	 	 else if (in == 3808) out = -298;
	 	 	 else if (in == 3809) out = -297;
	 	 	 else if (in == 3810) out = -296;
	 	 	 else if (in == 3811) out = -295;
	 	 	 else if (in == 3812) out = -294;
	 	 	 else if (in == 3813) out = -293;
	 	 	 else if (in == 3814) out = -292;
	 	 	 else if (in == 3815) out = -291;
	 	 	 else if (in == 3816) out = -290;
	 	 	 else if (in == 3817) out = -288;
	 	 	 else if (in == 3818) out = -287;
	 	 	 else if (in == 3819) out = -286;
	 	 	 else if (in == 3820) out = -285;
	 	 	 else if (in == 3821) out = -284;
	 	 	 else if (in == 3822) out = -283;
	 	 	 else if (in == 3823) out = -282;
	 	 	 else if (in == 3824) out = -281;
	 	 	 else if (in == 3825) out = -280;
	 	 	 else if (in == 3826) out = -279;
	 	 	 else if (in == 3827) out = -278;
	 	 	 else if (in == 3828) out = -277;
	 	 	 else if (in == 3829) out = -276;
	 	 	 else if (in == 3830) out = -275;
	 	 	 else if (in == 3831) out = -273;
	 	 	 else if (in == 3832) out = -272;
	 	 	 else if (in == 3833) out = -271;
	 	 	 else if (in == 3834) out = -270;
	 	 	 else if (in == 3835) out = -269;
	 	 	 else if (in == 3836) out = -268;
	 	 	 else if (in == 3837) out = -267;
	 	 	 else if (in == 3838) out = -266;
	 	 	 else if (in == 3839) out = -265;
	 	 	 else if (in == 3840) out = -264;
	 	 	 else if (in == 3841) out = -263;
	 	 	 else if (in == 3842) out = -262;
	 	 	 else if (in == 3843) out = -261;
	 	 	 else if (in == 3844) out = -260;
	 	 	 else if (in == 3845) out = -259;
	 	 	 else if (in == 3846) out = -257;
	 	 	 else if (in == 3847) out = -256;
	 	 	 else if (in == 3848) out = -255;
	 	 	 else if (in == 3849) out = -254;
	 	 	 else if (in == 3850) out = -253;
	 	 	 else if (in == 3851) out = -252;
	 	 	 else if (in == 3852) out = -251;
	 	 	 else if (in == 3853) out = -250;
	 	 	 else if (in == 3854) out = -249;
	 	 	 else if (in == 3855) out = -248;
	 	 	 else if (in == 3856) out = -247;
	 	 	 else if (in == 3857) out = -246;
	 	 	 else if (in == 3858) out = -245;
	 	 	 else if (in == 3859) out = -244;
	 	 	 else if (in == 3860) out = -243;
	 	 	 else if (in == 3861) out = -242;
	 	 	 else if (in == 3862) out = -240;
	 	 	 else if (in == 3863) out = -239;
	 	 	 else if (in == 3864) out = -238;
	 	 	 else if (in == 3865) out = -237;
	 	 	 else if (in == 3866) out = -236;
	 	 	 else if (in == 3867) out = -235;
	 	 	 else if (in == 3868) out = -234;
	 	 	 else if (in == 3869) out = -233;
	 	 	 else if (in == 3870) out = -232;
	 	 	 else if (in == 3871) out = -231;
	 	 	 else if (in == 3872) out = -230;
	 	 	 else if (in == 3873) out = -229;
	 	 	 else if (in == 3874) out = -228;
	 	 	 else if (in == 3875) out = -227;
	 	 	 else if (in == 3876) out = -226;
	 	 	 else if (in == 3877) out = -225;
	 	 	 else if (in == 3878) out = -224;
	 	 	 else if (in == 3879) out = -222;
	 	 	 else if (in == 3880) out = -221;
	 	 	 else if (in == 3881) out = -220;
	 	 	 else if (in == 3882) out = -219;
	 	 	 else if (in == 3883) out = -218;
	 	 	 else if (in == 3884) out = -217;
	 	 	 else if (in == 3885) out = -216;
	 	 	 else if (in == 3886) out = -215;
	 	 	 else if (in == 3887) out = -214;
	 	 	 else if (in == 3888) out = -213;
	 	 	 else if (in == 3889) out = -212;
	 	 	 else if (in == 3890) out = -211;
	 	 	 else if (in == 3891) out = -210;
	 	 	 else if (in == 3892) out = -209;
	 	 	 else if (in == 3893) out = -208;
	 	 	 else if (in == 3894) out = -207;
	 	 	 else if (in == 3895) out = -206;
	 	 	 else if (in == 3896) out = -205;
	 	 	 else if (in == 3897) out = -203;
	 	 	 else if (in == 3898) out = -202;
	 	 	 else if (in == 3899) out = -201;
	 	 	 else if (in == 3900) out = -200;
	 	 	 else if (in == 3901) out = -199;
	 	 	 else if (in == 3902) out = -198;
	 	 	 else if (in == 3903) out = -197;
	 	 	 else if (in == 3904) out = -196;
	 	 	 else if (in == 3905) out = -195;
	 	 	 else if (in == 3906) out = -194;
	 	 	 else if (in == 3907) out = -193;
	 	 	 else if (in == 3908) out = -192;
	 	 	 else if (in == 3909) out = -191;
	 	 	 else if (in == 3910) out = -190;
	 	 	 else if (in == 3911) out = -189;
	 	 	 else if (in == 3912) out = -188;
	 	 	 else if (in == 3913) out = -187;
	 	 	 else if (in == 3914) out = -186;
	 	 	 else if (in == 3915) out = -185;
	 	 	 else if (in == 3916) out = -184;
	 	 	 else if (in == 3917) out = -183;
	 	 	 else if (in == 3918) out = -181;
	 	 	 else if (in == 3919) out = -180;
	 	 	 else if (in == 3920) out = -179;
	 	 	 else if (in == 3921) out = -178;
	 	 	 else if (in == 3922) out = -177;
	 	 	 else if (in == 3923) out = -176;
	 	 	 else if (in == 3924) out = -175;
	 	 	 else if (in == 3925) out = -174;
	 	 	 else if (in == 3926) out = -173;
	 	 	 else if (in == 3927) out = -172;
	 	 	 else if (in == 3928) out = -171;
	 	 	 else if (in == 3929) out = -170;
	 	 	 else if (in == 3930) out = -169;
	 	 	 else if (in == 3931) out = -168;
	 	 	 else if (in == 3932) out = -167;
	 	 	 else if (in == 3933) out = -166;
	 	 	 else if (in == 3934) out = -165;
	 	 	 else if (in == 3935) out = -164;
	 	 	 else if (in == 3936) out = -163;
	 	 	 else if (in == 3937) out = -162;
	 	 	 else if (in == 3938) out = -161;
	 	 	 else if (in == 3939) out = -160;
	 	 	 else if (in == 3940) out = -159;
	 	 	 else if (in == 3941) out = -158;
	 	 	 else if (in == 3942) out = -156;
	 	 	 else if (in == 3943) out = -155;
	 	 	 else if (in == 3944) out = -154;
	 	 	 else if (in == 3945) out = -153;
	 	 	 else if (in == 3946) out = -152;
	 	 	 else if (in == 3947) out = -151;
	 	 	 else if (in == 3948) out = -150;
	 	 	 else if (in == 3949) out = -149;
	 	 	 else if (in == 3950) out = -148;
	 	 	 else if (in == 3951) out = -147;
	 	 	 else if (in == 3952) out = -146;
	 	 	 else if (in == 3953) out = -145;
	 	 	 else if (in == 3954) out = -144;
	 	 	 else if (in == 3955) out = -143;
	 	 	 else if (in == 3956) out = -142;
	 	 	 else if (in == 3957) out = -141;
	 	 	 else if (in == 3958) out = -140;
	 	 	 else if (in == 3959) out = -139;
	 	 	 else if (in == 3960) out = -138;
	 	 	 else if (in == 3961) out = -137;
	 	 	 else if (in == 3962) out = -136;
	 	 	 else if (in == 3963) out = -135;
	 	 	 else if (in == 3964) out = -134;
	 	 	 else if (in == 3965) out = -133;
	 	 	 else if (in == 3966) out = -132;
	 	 	 else if (in == 3967) out = -131;
	 	 	 else if (in == 3968) out = -130;
	 	 	 else if (in == 3969) out = -129;
	 	 	 else if (in == 3970) out = -127;
	 	 	 else if (in == 3971) out = -126;
	 	 	 else if (in == 3972) out = -125;
	 	 	 else if (in == 3973) out = -124;
	 	 	 else if (in == 3974) out = -123;
	 	 	 else if (in == 3975) out = -122;
	 	 	 else if (in == 3976) out = -121;
	 	 	 else if (in == 3977) out = -120;
	 	 	 else if (in == 3978) out = -119;
	 	 	 else if (in == 3979) out = -118;
	 	 	 else if (in == 3980) out = -117;
	 	 	 else if (in == 3981) out = -116;
	 	 	 else if (in == 3982) out = -115;
	 	 	 else if (in == 3983) out = -114;
	 	 	 else if (in == 3984) out = -113;
	 	 	 else if (in == 3985) out = -112;
	 	 	 else if (in == 3986) out = -111;
	 	 	 else if (in == 3987) out = -110;
	 	 	 else if (in == 3988) out = -109;
	 	 	 else if (in == 3989) out = -108;
	 	 	 else if (in == 3990) out = -107;
	 	 	 else if (in == 3991) out = -106;
	 	 	 else if (in == 3992) out = -105;
	 	 	 else if (in == 3993) out = -104;
	 	 	 else if (in == 3994) out = -103;
	 	 	 else if (in == 3995) out = -102;
	 	 	 else if (in == 3996) out = -101;
	 	 	 else if (in == 3997) out = -100;
	 	 	 else if (in == 3998) out = -99;
	 	 	 else if (in == 3999) out = -98;
	 	 	 else if (in == 4000) out = -97;
	 	 	 else if (in == 4001) out = -96;
	 	 	 else if (in == 4002) out = -95;
	 	 	 else if (in == 4003) out = -94;
	 	 	 else if (in == 4004) out = -93;
	 	 	 else if (in == 4005) out = -92;
	 	 	 else if (in == 4006) out = -91;
	 	 	 else if (in == 4007) out = -89;
	 	 	 else if (in == 4008) out = -88;
	 	 	 else if (in == 4009) out = -87;
	 	 	 else if (in == 4010) out = -86;
	 	 	 else if (in == 4011) out = -85;
	 	 	 else if (in == 4012) out = -84;
	 	 	 else if (in == 4013) out = -83;
	 	 	 else if (in == 4014) out = -82;
	 	 	 else if (in == 4015) out = -81;
	 	 	 else if (in == 4016) out = -80;
	 	 	 else if (in == 4017) out = -79;
	 	 	 else if (in == 4018) out = -78;
	 	 	 else if (in == 4019) out = -77;
	 	 	 else if (in == 4020) out = -76;
	 	 	 else if (in == 4021) out = -75;
	 	 	 else if (in == 4022) out = -74;
	 	 	 else if (in == 4023) out = -73;
	 	 	 else if (in == 4024) out = -72;
	 	 	 else if (in == 4025) out = -71;
	 	 	 else if (in == 4026) out = -70;
	 	 	 else if (in == 4027) out = -69;
	 	 	 else if (in == 4028) out = -68;
	 	 	 else if (in == 4029) out = -67;
	 	 	 else if (in == 4030) out = -66;
	 	 	 else if (in == 4031) out = -65;
	 	 	 else if (in == 4032) out = -64;
	 	 	 else if (in == 4033) out = -63;
	 	 	 else if (in == 4034) out = -62;
	 	 	 else if (in == 4035) out = -61;
	 	 	 else if (in == 4036) out = -60;
	 	 	 else if (in == 4037) out = -59;
	 	 	 else if (in == 4038) out = -58;
	 	 	 else if (in == 4039) out = -57;
	 	 	 else if (in == 4040) out = -56;
	 	 	 else if (in == 4041) out = -55;
	 	 	 else if (in == 4042) out = -54;
	 	 	 else if (in == 4043) out = -53;
	 	 	 else if (in == 4044) out = -52;
	 	 	 else if (in == 4045) out = -51;
	 	 	 else if (in == 4046) out = -50;
	 	 	 else if (in == 4047) out = -49;
	 	 	 else if (in == 4048) out = -48;
	 	 	 else if (in == 4049) out = -47;
	 	 	 else if (in == 4050) out = -46;
	 	 	 else if (in == 4051) out = -45;
	 	 	 else if (in == 4052) out = -44;
	 	 	 else if (in == 4053) out = -43;
	 	 	 else if (in == 4054) out = -42;
	 	 	 else if (in == 4055) out = -41;
	 	 	 else if (in == 4056) out = -40;
	 	 	 else if (in == 4057) out = -39;
	 	 	 else if (in == 4058) out = -38;
	 	 	 else if (in == 4059) out = -37;
	 	 	 else if (in == 4060) out = -36;
	 	 	 else if (in == 4061) out = -35;
	 	 	 else if (in == 4062) out = -34;
	 	 	 else if (in == 4063) out = -33;
	 	 	 else if (in == 4064) out = -32;
	 	 	 else if (in == 4065) out = -31;
	 	 	 else if (in == 4066) out = -30;
	 	 	 else if (in == 4067) out = -29;
	 	 	 else if (in == 4068) out = -28;
	 	 	 else if (in == 4069) out = -27;
	 	 	 else if (in == 4070) out = -26;
	 	 	 else if (in == 4071) out = -25;
	 	 	 else if (in == 4072) out = -24;
	 	 	 else if (in == 4073) out = -23;
	 	 	 else if (in == 4074) out = -22;
	 	 	 else if (in == 4075) out = -21;
	 	 	 else if (in == 4076) out = -20;
	 	 	 else if (in == 4077) out = -19;
	 	 	 else if (in == 4078) out = -18;
	 	 	 else if (in == 4079) out = -17;
	 	 	 else if (in == 4080) out = -16;
	 	 	 else if (in == 4081) out = -15;
	 	 	 else if (in == 4082) out = -14;
	 	 	 else if (in == 4083) out = -13;
	 	 	 else if (in == 4084) out = -12;
	 	 	 else if (in == 4085) out = -11;
	 	 	 else if (in == 4086) out = -10;
	 	 	 else if (in == 4087) out = -9;
	 	 	 else if (in == 4088) out = -8;
	 	 	 else if (in == 4089) out = -7;
	 	 	 else if (in == 4090) out = -6;
	 	 	 else if (in == 4091) out = -5;
	 	 	 else if (in == 4092) out = -4;
	 	 	 else if (in == 4093) out = -3;
	 	 	 else if (in == 4094) out = -2;
	 	 	 else if (in == 4095) out = -1;
	 	 	 else if (in == 4096) out = 0;
	 	 	else out=0;
	 endmodule