`ifndef header
`define header
    parameter ROWS = 1; // Number of Rows
    parameter COLUMNS = 2; // Number of Columns
`endif
